`timescale 1ns / 1ps

module MinSADFinder(SADValues, MinI, MinJ, MinVal);

    input [64*64*12-1:0] SADValues;
    output wire [5:0] MinI, MinJ;
    output wire [11:0] MinVal;

    wire [11:0] comp0minVal;
    wire [5:0] comp0minI, comp0minJ;
    Comparator comp0(SADValues[0*12 +: 12], 0, 0, SADValues[0*12 +: 12], 0, 0, comp0minVal, comp0minI, comp0minJ);
    wire [11:0] comp1minVal;
    wire [5:0] comp1minI, comp1minJ;
    Comparator comp1(SADValues[1*12 +: 12], 0, 1, SADValues[64*12 +: 12], 1, 0, comp1minVal, comp1minI, comp1minJ);
    wire [11:0] comp2minVal;
    wire [5:0] comp2minI, comp2minJ;
    Comparator comp2(SADValues[128*12 +: 12], 2, 0, SADValues[65*12 +: 12], 1, 1, comp2minVal, comp2minI, comp2minJ);
    wire [11:0] comp3minVal;
    wire [5:0] comp3minI, comp3minJ;
    Comparator comp3(SADValues[2*12 +: 12], 0, 2, SADValues[3*12 +: 12], 0, 3, comp3minVal, comp3minI, comp3minJ);
    wire [11:0] comp4minVal;
    wire [5:0] comp4minI, comp4minJ;
    Comparator comp4(SADValues[66*12 +: 12], 1, 2, SADValues[129*12 +: 12], 2, 1, comp4minVal, comp4minI, comp4minJ);
    wire [11:0] comp5minVal;
    wire [5:0] comp5minI, comp5minJ;
    Comparator comp5(SADValues[192*12 +: 12], 3, 0, SADValues[256*12 +: 12], 4, 0, comp5minVal, comp5minI, comp5minJ);
    wire [11:0] comp6minVal;
    wire [5:0] comp6minI, comp6minJ;
    Comparator comp6(SADValues[193*12 +: 12], 3, 1, SADValues[130*12 +: 12], 2, 2, comp6minVal, comp6minI, comp6minJ);
    wire [11:0] comp7minVal;
    wire [5:0] comp7minI, comp7minJ;
    Comparator comp7(SADValues[67*12 +: 12], 1, 3, SADValues[4*12 +: 12], 0, 4, comp7minVal, comp7minI, comp7minJ);
    wire [11:0] comp8minVal;
    wire [5:0] comp8minI, comp8minJ;
    Comparator comp8(SADValues[5*12 +: 12], 0, 5, SADValues[68*12 +: 12], 1, 4, comp8minVal, comp8minI, comp8minJ);
    wire [11:0] comp9minVal;
    wire [5:0] comp9minI, comp9minJ;
    Comparator comp9(SADValues[131*12 +: 12], 2, 3, SADValues[194*12 +: 12], 3, 2, comp9minVal, comp9minI, comp9minJ);
    wire [11:0] comp10minVal;
    wire [5:0] comp10minI, comp10minJ;
    Comparator comp10(SADValues[257*12 +: 12], 4, 1, SADValues[320*12 +: 12], 5, 0, comp10minVal, comp10minI, comp10minJ);
    wire [11:0] comp11minVal;
    wire [5:0] comp11minI, comp11minJ;
    Comparator comp11(SADValues[384*12 +: 12], 6, 0, SADValues[321*12 +: 12], 5, 1, comp11minVal, comp11minI, comp11minJ);
    wire [11:0] comp12minVal;
    wire [5:0] comp12minI, comp12minJ;
    Comparator comp12(SADValues[258*12 +: 12], 4, 2, SADValues[195*12 +: 12], 3, 3, comp12minVal, comp12minI, comp12minJ);
    wire [11:0] comp13minVal;
    wire [5:0] comp13minI, comp13minJ;
    Comparator comp13(SADValues[132*12 +: 12], 2, 4, SADValues[69*12 +: 12], 1, 5, comp13minVal, comp13minI, comp13minJ);
    wire [11:0] comp14minVal;
    wire [5:0] comp14minI, comp14minJ;
    Comparator comp14(SADValues[6*12 +: 12], 0, 6, SADValues[7*12 +: 12], 0, 7, comp14minVal, comp14minI, comp14minJ);
    wire [11:0] comp15minVal;
    wire [5:0] comp15minI, comp15minJ;
    Comparator comp15(SADValues[70*12 +: 12], 1, 6, SADValues[133*12 +: 12], 2, 5, comp15minVal, comp15minI, comp15minJ);
    wire [11:0] comp16minVal;
    wire [5:0] comp16minI, comp16minJ;
    Comparator comp16(SADValues[196*12 +: 12], 3, 4, SADValues[259*12 +: 12], 4, 3, comp16minVal, comp16minI, comp16minJ);
    wire [11:0] comp17minVal;
    wire [5:0] comp17minI, comp17minJ;
    Comparator comp17(SADValues[322*12 +: 12], 5, 2, SADValues[385*12 +: 12], 6, 1, comp17minVal, comp17minI, comp17minJ);
    wire [11:0] comp18minVal;
    wire [5:0] comp18minI, comp18minJ;
    Comparator comp18(SADValues[448*12 +: 12], 7, 0, SADValues[512*12 +: 12], 8, 0, comp18minVal, comp18minI, comp18minJ);
    wire [11:0] comp19minVal;
    wire [5:0] comp19minI, comp19minJ;
    Comparator comp19(SADValues[449*12 +: 12], 7, 1, SADValues[386*12 +: 12], 6, 2, comp19minVal, comp19minI, comp19minJ);
    wire [11:0] comp20minVal;
    wire [5:0] comp20minI, comp20minJ;
    Comparator comp20(SADValues[323*12 +: 12], 5, 3, SADValues[260*12 +: 12], 4, 4, comp20minVal, comp20minI, comp20minJ);
    wire [11:0] comp21minVal;
    wire [5:0] comp21minI, comp21minJ;
    Comparator comp21(SADValues[197*12 +: 12], 3, 5, SADValues[134*12 +: 12], 2, 6, comp21minVal, comp21minI, comp21minJ);
    wire [11:0] comp22minVal;
    wire [5:0] comp22minI, comp22minJ;
    Comparator comp22(SADValues[71*12 +: 12], 1, 7, SADValues[8*12 +: 12], 0, 8, comp22minVal, comp22minI, comp22minJ);
    wire [11:0] comp23minVal;
    wire [5:0] comp23minI, comp23minJ;
    Comparator comp23(SADValues[9*12 +: 12], 0, 9, SADValues[72*12 +: 12], 1, 8, comp23minVal, comp23minI, comp23minJ);
    wire [11:0] comp24minVal;
    wire [5:0] comp24minI, comp24minJ;
    Comparator comp24(SADValues[135*12 +: 12], 2, 7, SADValues[198*12 +: 12], 3, 6, comp24minVal, comp24minI, comp24minJ);
    wire [11:0] comp25minVal;
    wire [5:0] comp25minI, comp25minJ;
    Comparator comp25(SADValues[261*12 +: 12], 4, 5, SADValues[324*12 +: 12], 5, 4, comp25minVal, comp25minI, comp25minJ);
    wire [11:0] comp26minVal;
    wire [5:0] comp26minI, comp26minJ;
    Comparator comp26(SADValues[387*12 +: 12], 6, 3, SADValues[450*12 +: 12], 7, 2, comp26minVal, comp26minI, comp26minJ);
    wire [11:0] comp27minVal;
    wire [5:0] comp27minI, comp27minJ;
    Comparator comp27(SADValues[513*12 +: 12], 8, 1, SADValues[576*12 +: 12], 9, 0, comp27minVal, comp27minI, comp27minJ);
    wire [11:0] comp28minVal;
    wire [5:0] comp28minI, comp28minJ;
    Comparator comp28(SADValues[640*12 +: 12], 10, 0, SADValues[577*12 +: 12], 9, 1, comp28minVal, comp28minI, comp28minJ);
    wire [11:0] comp29minVal;
    wire [5:0] comp29minI, comp29minJ;
    Comparator comp29(SADValues[514*12 +: 12], 8, 2, SADValues[451*12 +: 12], 7, 3, comp29minVal, comp29minI, comp29minJ);
    wire [11:0] comp30minVal;
    wire [5:0] comp30minI, comp30minJ;
    Comparator comp30(SADValues[388*12 +: 12], 6, 4, SADValues[325*12 +: 12], 5, 5, comp30minVal, comp30minI, comp30minJ);
    wire [11:0] comp31minVal;
    wire [5:0] comp31minI, comp31minJ;
    Comparator comp31(SADValues[262*12 +: 12], 4, 6, SADValues[199*12 +: 12], 3, 7, comp31minVal, comp31minI, comp31minJ);
    wire [11:0] comp32minVal;
    wire [5:0] comp32minI, comp32minJ;
    Comparator comp32(SADValues[136*12 +: 12], 2, 8, SADValues[73*12 +: 12], 1, 9, comp32minVal, comp32minI, comp32minJ);
    wire [11:0] comp33minVal;
    wire [5:0] comp33minI, comp33minJ;
    Comparator comp33(SADValues[10*12 +: 12], 0, 10, SADValues[11*12 +: 12], 0, 11, comp33minVal, comp33minI, comp33minJ);
    wire [11:0] comp34minVal;
    wire [5:0] comp34minI, comp34minJ;
    Comparator comp34(SADValues[74*12 +: 12], 1, 10, SADValues[137*12 +: 12], 2, 9, comp34minVal, comp34minI, comp34minJ);
    wire [11:0] comp35minVal;
    wire [5:0] comp35minI, comp35minJ;
    Comparator comp35(SADValues[200*12 +: 12], 3, 8, SADValues[263*12 +: 12], 4, 7, comp35minVal, comp35minI, comp35minJ);
    wire [11:0] comp36minVal;
    wire [5:0] comp36minI, comp36minJ;
    Comparator comp36(SADValues[326*12 +: 12], 5, 6, SADValues[389*12 +: 12], 6, 5, comp36minVal, comp36minI, comp36minJ);
    wire [11:0] comp37minVal;
    wire [5:0] comp37minI, comp37minJ;
    Comparator comp37(SADValues[452*12 +: 12], 7, 4, SADValues[515*12 +: 12], 8, 3, comp37minVal, comp37minI, comp37minJ);
    wire [11:0] comp38minVal;
    wire [5:0] comp38minI, comp38minJ;
    Comparator comp38(SADValues[578*12 +: 12], 9, 2, SADValues[641*12 +: 12], 10, 1, comp38minVal, comp38minI, comp38minJ);
    wire [11:0] comp39minVal;
    wire [5:0] comp39minI, comp39minJ;
    Comparator comp39(SADValues[704*12 +: 12], 11, 0, SADValues[768*12 +: 12], 12, 0, comp39minVal, comp39minI, comp39minJ);
    wire [11:0] comp40minVal;
    wire [5:0] comp40minI, comp40minJ;
    Comparator comp40(SADValues[705*12 +: 12], 11, 1, SADValues[642*12 +: 12], 10, 2, comp40minVal, comp40minI, comp40minJ);
    wire [11:0] comp41minVal;
    wire [5:0] comp41minI, comp41minJ;
    Comparator comp41(SADValues[579*12 +: 12], 9, 3, SADValues[516*12 +: 12], 8, 4, comp41minVal, comp41minI, comp41minJ);
    wire [11:0] comp42minVal;
    wire [5:0] comp42minI, comp42minJ;
    Comparator comp42(SADValues[453*12 +: 12], 7, 5, SADValues[390*12 +: 12], 6, 6, comp42minVal, comp42minI, comp42minJ);
    wire [11:0] comp43minVal;
    wire [5:0] comp43minI, comp43minJ;
    Comparator comp43(SADValues[327*12 +: 12], 5, 7, SADValues[264*12 +: 12], 4, 8, comp43minVal, comp43minI, comp43minJ);
    wire [11:0] comp44minVal;
    wire [5:0] comp44minI, comp44minJ;
    Comparator comp44(SADValues[201*12 +: 12], 3, 9, SADValues[138*12 +: 12], 2, 10, comp44minVal, comp44minI, comp44minJ);
    wire [11:0] comp45minVal;
    wire [5:0] comp45minI, comp45minJ;
    Comparator comp45(SADValues[75*12 +: 12], 1, 11, SADValues[12*12 +: 12], 0, 12, comp45minVal, comp45minI, comp45minJ);
    wire [11:0] comp46minVal;
    wire [5:0] comp46minI, comp46minJ;
    Comparator comp46(SADValues[13*12 +: 12], 0, 13, SADValues[76*12 +: 12], 1, 12, comp46minVal, comp46minI, comp46minJ);
    wire [11:0] comp47minVal;
    wire [5:0] comp47minI, comp47minJ;
    Comparator comp47(SADValues[139*12 +: 12], 2, 11, SADValues[202*12 +: 12], 3, 10, comp47minVal, comp47minI, comp47minJ);
    wire [11:0] comp48minVal;
    wire [5:0] comp48minI, comp48minJ;
    Comparator comp48(SADValues[265*12 +: 12], 4, 9, SADValues[328*12 +: 12], 5, 8, comp48minVal, comp48minI, comp48minJ);
    wire [11:0] comp49minVal;
    wire [5:0] comp49minI, comp49minJ;
    Comparator comp49(SADValues[391*12 +: 12], 6, 7, SADValues[454*12 +: 12], 7, 6, comp49minVal, comp49minI, comp49minJ);
    wire [11:0] comp50minVal;
    wire [5:0] comp50minI, comp50minJ;
    Comparator comp50(SADValues[517*12 +: 12], 8, 5, SADValues[580*12 +: 12], 9, 4, comp50minVal, comp50minI, comp50minJ);
    wire [11:0] comp51minVal;
    wire [5:0] comp51minI, comp51minJ;
    Comparator comp51(SADValues[643*12 +: 12], 10, 3, SADValues[706*12 +: 12], 11, 2, comp51minVal, comp51minI, comp51minJ);
    wire [11:0] comp52minVal;
    wire [5:0] comp52minI, comp52minJ;
    Comparator comp52(SADValues[769*12 +: 12], 12, 1, SADValues[832*12 +: 12], 13, 0, comp52minVal, comp52minI, comp52minJ);
    wire [11:0] comp53minVal;
    wire [5:0] comp53minI, comp53minJ;
    Comparator comp53(SADValues[896*12 +: 12], 14, 0, SADValues[833*12 +: 12], 13, 1, comp53minVal, comp53minI, comp53minJ);
    wire [11:0] comp54minVal;
    wire [5:0] comp54minI, comp54minJ;
    Comparator comp54(SADValues[770*12 +: 12], 12, 2, SADValues[707*12 +: 12], 11, 3, comp54minVal, comp54minI, comp54minJ);
    wire [11:0] comp55minVal;
    wire [5:0] comp55minI, comp55minJ;
    Comparator comp55(SADValues[644*12 +: 12], 10, 4, SADValues[581*12 +: 12], 9, 5, comp55minVal, comp55minI, comp55minJ);
    wire [11:0] comp56minVal;
    wire [5:0] comp56minI, comp56minJ;
    Comparator comp56(SADValues[518*12 +: 12], 8, 6, SADValues[455*12 +: 12], 7, 7, comp56minVal, comp56minI, comp56minJ);
    wire [11:0] comp57minVal;
    wire [5:0] comp57minI, comp57minJ;
    Comparator comp57(SADValues[392*12 +: 12], 6, 8, SADValues[329*12 +: 12], 5, 9, comp57minVal, comp57minI, comp57minJ);
    wire [11:0] comp58minVal;
    wire [5:0] comp58minI, comp58minJ;
    Comparator comp58(SADValues[266*12 +: 12], 4, 10, SADValues[203*12 +: 12], 3, 11, comp58minVal, comp58minI, comp58minJ);
    wire [11:0] comp59minVal;
    wire [5:0] comp59minI, comp59minJ;
    Comparator comp59(SADValues[140*12 +: 12], 2, 12, SADValues[77*12 +: 12], 1, 13, comp59minVal, comp59minI, comp59minJ);
    wire [11:0] comp60minVal;
    wire [5:0] comp60minI, comp60minJ;
    Comparator comp60(SADValues[14*12 +: 12], 0, 14, SADValues[15*12 +: 12], 0, 15, comp60minVal, comp60minI, comp60minJ);
    wire [11:0] comp61minVal;
    wire [5:0] comp61minI, comp61minJ;
    Comparator comp61(SADValues[78*12 +: 12], 1, 14, SADValues[141*12 +: 12], 2, 13, comp61minVal, comp61minI, comp61minJ);
    wire [11:0] comp62minVal;
    wire [5:0] comp62minI, comp62minJ;
    Comparator comp62(SADValues[204*12 +: 12], 3, 12, SADValues[267*12 +: 12], 4, 11, comp62minVal, comp62minI, comp62minJ);
    wire [11:0] comp63minVal;
    wire [5:0] comp63minI, comp63minJ;
    Comparator comp63(SADValues[330*12 +: 12], 5, 10, SADValues[393*12 +: 12], 6, 9, comp63minVal, comp63minI, comp63minJ);
    wire [11:0] comp64minVal;
    wire [5:0] comp64minI, comp64minJ;
    Comparator comp64(SADValues[456*12 +: 12], 7, 8, SADValues[519*12 +: 12], 8, 7, comp64minVal, comp64minI, comp64minJ);
    wire [11:0] comp65minVal;
    wire [5:0] comp65minI, comp65minJ;
    Comparator comp65(SADValues[582*12 +: 12], 9, 6, SADValues[645*12 +: 12], 10, 5, comp65minVal, comp65minI, comp65minJ);
    wire [11:0] comp66minVal;
    wire [5:0] comp66minI, comp66minJ;
    Comparator comp66(SADValues[708*12 +: 12], 11, 4, SADValues[771*12 +: 12], 12, 3, comp66minVal, comp66minI, comp66minJ);
    wire [11:0] comp67minVal;
    wire [5:0] comp67minI, comp67minJ;
    Comparator comp67(SADValues[834*12 +: 12], 13, 2, SADValues[897*12 +: 12], 14, 1, comp67minVal, comp67minI, comp67minJ);
    wire [11:0] comp68minVal;
    wire [5:0] comp68minI, comp68minJ;
    Comparator comp68(SADValues[960*12 +: 12], 15, 0, SADValues[1024*12 +: 12], 16, 0, comp68minVal, comp68minI, comp68minJ);
    wire [11:0] comp69minVal;
    wire [5:0] comp69minI, comp69minJ;
    Comparator comp69(SADValues[961*12 +: 12], 15, 1, SADValues[898*12 +: 12], 14, 2, comp69minVal, comp69minI, comp69minJ);
    wire [11:0] comp70minVal;
    wire [5:0] comp70minI, comp70minJ;
    Comparator comp70(SADValues[835*12 +: 12], 13, 3, SADValues[772*12 +: 12], 12, 4, comp70minVal, comp70minI, comp70minJ);
    wire [11:0] comp71minVal;
    wire [5:0] comp71minI, comp71minJ;
    Comparator comp71(SADValues[709*12 +: 12], 11, 5, SADValues[646*12 +: 12], 10, 6, comp71minVal, comp71minI, comp71minJ);
    wire [11:0] comp72minVal;
    wire [5:0] comp72minI, comp72minJ;
    Comparator comp72(SADValues[583*12 +: 12], 9, 7, SADValues[520*12 +: 12], 8, 8, comp72minVal, comp72minI, comp72minJ);
    wire [11:0] comp73minVal;
    wire [5:0] comp73minI, comp73minJ;
    Comparator comp73(SADValues[457*12 +: 12], 7, 9, SADValues[394*12 +: 12], 6, 10, comp73minVal, comp73minI, comp73minJ);
    wire [11:0] comp74minVal;
    wire [5:0] comp74minI, comp74minJ;
    Comparator comp74(SADValues[331*12 +: 12], 5, 11, SADValues[268*12 +: 12], 4, 12, comp74minVal, comp74minI, comp74minJ);
    wire [11:0] comp75minVal;
    wire [5:0] comp75minI, comp75minJ;
    Comparator comp75(SADValues[205*12 +: 12], 3, 13, SADValues[142*12 +: 12], 2, 14, comp75minVal, comp75minI, comp75minJ);
    wire [11:0] comp76minVal;
    wire [5:0] comp76minI, comp76minJ;
    Comparator comp76(SADValues[79*12 +: 12], 1, 15, SADValues[16*12 +: 12], 0, 16, comp76minVal, comp76minI, comp76minJ);
    wire [11:0] comp77minVal;
    wire [5:0] comp77minI, comp77minJ;
    Comparator comp77(SADValues[17*12 +: 12], 0, 17, SADValues[80*12 +: 12], 1, 16, comp77minVal, comp77minI, comp77minJ);
    wire [11:0] comp78minVal;
    wire [5:0] comp78minI, comp78minJ;
    Comparator comp78(SADValues[143*12 +: 12], 2, 15, SADValues[206*12 +: 12], 3, 14, comp78minVal, comp78minI, comp78minJ);
    wire [11:0] comp79minVal;
    wire [5:0] comp79minI, comp79minJ;
    Comparator comp79(SADValues[269*12 +: 12], 4, 13, SADValues[332*12 +: 12], 5, 12, comp79minVal, comp79minI, comp79minJ);
    wire [11:0] comp80minVal;
    wire [5:0] comp80minI, comp80minJ;
    Comparator comp80(SADValues[395*12 +: 12], 6, 11, SADValues[458*12 +: 12], 7, 10, comp80minVal, comp80minI, comp80minJ);
    wire [11:0] comp81minVal;
    wire [5:0] comp81minI, comp81minJ;
    Comparator comp81(SADValues[521*12 +: 12], 8, 9, SADValues[584*12 +: 12], 9, 8, comp81minVal, comp81minI, comp81minJ);
    wire [11:0] comp82minVal;
    wire [5:0] comp82minI, comp82minJ;
    Comparator comp82(SADValues[647*12 +: 12], 10, 7, SADValues[710*12 +: 12], 11, 6, comp82minVal, comp82minI, comp82minJ);
    wire [11:0] comp83minVal;
    wire [5:0] comp83minI, comp83minJ;
    Comparator comp83(SADValues[773*12 +: 12], 12, 5, SADValues[836*12 +: 12], 13, 4, comp83minVal, comp83minI, comp83minJ);
    wire [11:0] comp84minVal;
    wire [5:0] comp84minI, comp84minJ;
    Comparator comp84(SADValues[899*12 +: 12], 14, 3, SADValues[962*12 +: 12], 15, 2, comp84minVal, comp84minI, comp84minJ);
    wire [11:0] comp85minVal;
    wire [5:0] comp85minI, comp85minJ;
    Comparator comp85(SADValues[1025*12 +: 12], 16, 1, SADValues[1088*12 +: 12], 17, 0, comp85minVal, comp85minI, comp85minJ);
    wire [11:0] comp86minVal;
    wire [5:0] comp86minI, comp86minJ;
    Comparator comp86(SADValues[1152*12 +: 12], 18, 0, SADValues[1089*12 +: 12], 17, 1, comp86minVal, comp86minI, comp86minJ);
    wire [11:0] comp87minVal;
    wire [5:0] comp87minI, comp87minJ;
    Comparator comp87(SADValues[1026*12 +: 12], 16, 2, SADValues[963*12 +: 12], 15, 3, comp87minVal, comp87minI, comp87minJ);
    wire [11:0] comp88minVal;
    wire [5:0] comp88minI, comp88minJ;
    Comparator comp88(SADValues[900*12 +: 12], 14, 4, SADValues[837*12 +: 12], 13, 5, comp88minVal, comp88minI, comp88minJ);
    wire [11:0] comp89minVal;
    wire [5:0] comp89minI, comp89minJ;
    Comparator comp89(SADValues[774*12 +: 12], 12, 6, SADValues[711*12 +: 12], 11, 7, comp89minVal, comp89minI, comp89minJ);
    wire [11:0] comp90minVal;
    wire [5:0] comp90minI, comp90minJ;
    Comparator comp90(SADValues[648*12 +: 12], 10, 8, SADValues[585*12 +: 12], 9, 9, comp90minVal, comp90minI, comp90minJ);
    wire [11:0] comp91minVal;
    wire [5:0] comp91minI, comp91minJ;
    Comparator comp91(SADValues[522*12 +: 12], 8, 10, SADValues[459*12 +: 12], 7, 11, comp91minVal, comp91minI, comp91minJ);
    wire [11:0] comp92minVal;
    wire [5:0] comp92minI, comp92minJ;
    Comparator comp92(SADValues[396*12 +: 12], 6, 12, SADValues[333*12 +: 12], 5, 13, comp92minVal, comp92minI, comp92minJ);
    wire [11:0] comp93minVal;
    wire [5:0] comp93minI, comp93minJ;
    Comparator comp93(SADValues[270*12 +: 12], 4, 14, SADValues[207*12 +: 12], 3, 15, comp93minVal, comp93minI, comp93minJ);
    wire [11:0] comp94minVal;
    wire [5:0] comp94minI, comp94minJ;
    Comparator comp94(SADValues[144*12 +: 12], 2, 16, SADValues[81*12 +: 12], 1, 17, comp94minVal, comp94minI, comp94minJ);
    wire [11:0] comp95minVal;
    wire [5:0] comp95minI, comp95minJ;
    Comparator comp95(SADValues[18*12 +: 12], 0, 18, SADValues[19*12 +: 12], 0, 19, comp95minVal, comp95minI, comp95minJ);
    wire [11:0] comp96minVal;
    wire [5:0] comp96minI, comp96minJ;
    Comparator comp96(SADValues[82*12 +: 12], 1, 18, SADValues[145*12 +: 12], 2, 17, comp96minVal, comp96minI, comp96minJ);
    wire [11:0] comp97minVal;
    wire [5:0] comp97minI, comp97minJ;
    Comparator comp97(SADValues[208*12 +: 12], 3, 16, SADValues[271*12 +: 12], 4, 15, comp97minVal, comp97minI, comp97minJ);
    wire [11:0] comp98minVal;
    wire [5:0] comp98minI, comp98minJ;
    Comparator comp98(SADValues[334*12 +: 12], 5, 14, SADValues[397*12 +: 12], 6, 13, comp98minVal, comp98minI, comp98minJ);
    wire [11:0] comp99minVal;
    wire [5:0] comp99minI, comp99minJ;
    Comparator comp99(SADValues[460*12 +: 12], 7, 12, SADValues[523*12 +: 12], 8, 11, comp99minVal, comp99minI, comp99minJ);
    wire [11:0] comp100minVal;
    wire [5:0] comp100minI, comp100minJ;
    Comparator comp100(SADValues[586*12 +: 12], 9, 10, SADValues[649*12 +: 12], 10, 9, comp100minVal, comp100minI, comp100minJ);
    wire [11:0] comp101minVal;
    wire [5:0] comp101minI, comp101minJ;
    Comparator comp101(SADValues[712*12 +: 12], 11, 8, SADValues[775*12 +: 12], 12, 7, comp101minVal, comp101minI, comp101minJ);
    wire [11:0] comp102minVal;
    wire [5:0] comp102minI, comp102minJ;
    Comparator comp102(SADValues[838*12 +: 12], 13, 6, SADValues[901*12 +: 12], 14, 5, comp102minVal, comp102minI, comp102minJ);
    wire [11:0] comp103minVal;
    wire [5:0] comp103minI, comp103minJ;
    Comparator comp103(SADValues[964*12 +: 12], 15, 4, SADValues[1027*12 +: 12], 16, 3, comp103minVal, comp103minI, comp103minJ);
    wire [11:0] comp104minVal;
    wire [5:0] comp104minI, comp104minJ;
    Comparator comp104(SADValues[1090*12 +: 12], 17, 2, SADValues[1153*12 +: 12], 18, 1, comp104minVal, comp104minI, comp104minJ);
    wire [11:0] comp105minVal;
    wire [5:0] comp105minI, comp105minJ;
    Comparator comp105(SADValues[1216*12 +: 12], 19, 0, SADValues[1280*12 +: 12], 20, 0, comp105minVal, comp105minI, comp105minJ);
    wire [11:0] comp106minVal;
    wire [5:0] comp106minI, comp106minJ;
    Comparator comp106(SADValues[1217*12 +: 12], 19, 1, SADValues[1154*12 +: 12], 18, 2, comp106minVal, comp106minI, comp106minJ);
    wire [11:0] comp107minVal;
    wire [5:0] comp107minI, comp107minJ;
    Comparator comp107(SADValues[1091*12 +: 12], 17, 3, SADValues[1028*12 +: 12], 16, 4, comp107minVal, comp107minI, comp107minJ);
    wire [11:0] comp108minVal;
    wire [5:0] comp108minI, comp108minJ;
    Comparator comp108(SADValues[965*12 +: 12], 15, 5, SADValues[902*12 +: 12], 14, 6, comp108minVal, comp108minI, comp108minJ);
    wire [11:0] comp109minVal;
    wire [5:0] comp109minI, comp109minJ;
    Comparator comp109(SADValues[839*12 +: 12], 13, 7, SADValues[776*12 +: 12], 12, 8, comp109minVal, comp109minI, comp109minJ);
    wire [11:0] comp110minVal;
    wire [5:0] comp110minI, comp110minJ;
    Comparator comp110(SADValues[713*12 +: 12], 11, 9, SADValues[650*12 +: 12], 10, 10, comp110minVal, comp110minI, comp110minJ);
    wire [11:0] comp111minVal;
    wire [5:0] comp111minI, comp111minJ;
    Comparator comp111(SADValues[587*12 +: 12], 9, 11, SADValues[524*12 +: 12], 8, 12, comp111minVal, comp111minI, comp111minJ);
    wire [11:0] comp112minVal;
    wire [5:0] comp112minI, comp112minJ;
    Comparator comp112(SADValues[461*12 +: 12], 7, 13, SADValues[398*12 +: 12], 6, 14, comp112minVal, comp112minI, comp112minJ);
    wire [11:0] comp113minVal;
    wire [5:0] comp113minI, comp113minJ;
    Comparator comp113(SADValues[335*12 +: 12], 5, 15, SADValues[272*12 +: 12], 4, 16, comp113minVal, comp113minI, comp113minJ);
    wire [11:0] comp114minVal;
    wire [5:0] comp114minI, comp114minJ;
    Comparator comp114(SADValues[209*12 +: 12], 3, 17, SADValues[146*12 +: 12], 2, 18, comp114minVal, comp114minI, comp114minJ);
    wire [11:0] comp115minVal;
    wire [5:0] comp115minI, comp115minJ;
    Comparator comp115(SADValues[83*12 +: 12], 1, 19, SADValues[20*12 +: 12], 0, 20, comp115minVal, comp115minI, comp115minJ);
    wire [11:0] comp116minVal;
    wire [5:0] comp116minI, comp116minJ;
    Comparator comp116(SADValues[21*12 +: 12], 0, 21, SADValues[84*12 +: 12], 1, 20, comp116minVal, comp116minI, comp116minJ);
    wire [11:0] comp117minVal;
    wire [5:0] comp117minI, comp117minJ;
    Comparator comp117(SADValues[147*12 +: 12], 2, 19, SADValues[210*12 +: 12], 3, 18, comp117minVal, comp117minI, comp117minJ);
    wire [11:0] comp118minVal;
    wire [5:0] comp118minI, comp118minJ;
    Comparator comp118(SADValues[273*12 +: 12], 4, 17, SADValues[336*12 +: 12], 5, 16, comp118minVal, comp118minI, comp118minJ);
    wire [11:0] comp119minVal;
    wire [5:0] comp119minI, comp119minJ;
    Comparator comp119(SADValues[399*12 +: 12], 6, 15, SADValues[462*12 +: 12], 7, 14, comp119minVal, comp119minI, comp119minJ);
    wire [11:0] comp120minVal;
    wire [5:0] comp120minI, comp120minJ;
    Comparator comp120(SADValues[525*12 +: 12], 8, 13, SADValues[588*12 +: 12], 9, 12, comp120minVal, comp120minI, comp120minJ);
    wire [11:0] comp121minVal;
    wire [5:0] comp121minI, comp121minJ;
    Comparator comp121(SADValues[651*12 +: 12], 10, 11, SADValues[714*12 +: 12], 11, 10, comp121minVal, comp121minI, comp121minJ);
    wire [11:0] comp122minVal;
    wire [5:0] comp122minI, comp122minJ;
    Comparator comp122(SADValues[777*12 +: 12], 12, 9, SADValues[840*12 +: 12], 13, 8, comp122minVal, comp122minI, comp122minJ);
    wire [11:0] comp123minVal;
    wire [5:0] comp123minI, comp123minJ;
    Comparator comp123(SADValues[903*12 +: 12], 14, 7, SADValues[966*12 +: 12], 15, 6, comp123minVal, comp123minI, comp123minJ);
    wire [11:0] comp124minVal;
    wire [5:0] comp124minI, comp124minJ;
    Comparator comp124(SADValues[1029*12 +: 12], 16, 5, SADValues[1092*12 +: 12], 17, 4, comp124minVal, comp124minI, comp124minJ);
    wire [11:0] comp125minVal;
    wire [5:0] comp125minI, comp125minJ;
    Comparator comp125(SADValues[1155*12 +: 12], 18, 3, SADValues[1218*12 +: 12], 19, 2, comp125minVal, comp125minI, comp125minJ);
    wire [11:0] comp126minVal;
    wire [5:0] comp126minI, comp126minJ;
    Comparator comp126(SADValues[1281*12 +: 12], 20, 1, SADValues[1344*12 +: 12], 21, 0, comp126minVal, comp126minI, comp126minJ);
    wire [11:0] comp127minVal;
    wire [5:0] comp127minI, comp127minJ;
    Comparator comp127(SADValues[1408*12 +: 12], 22, 0, SADValues[1345*12 +: 12], 21, 1, comp127minVal, comp127minI, comp127minJ);
    wire [11:0] comp128minVal;
    wire [5:0] comp128minI, comp128minJ;
    Comparator comp128(SADValues[1282*12 +: 12], 20, 2, SADValues[1219*12 +: 12], 19, 3, comp128minVal, comp128minI, comp128minJ);
    wire [11:0] comp129minVal;
    wire [5:0] comp129minI, comp129minJ;
    Comparator comp129(SADValues[1156*12 +: 12], 18, 4, SADValues[1093*12 +: 12], 17, 5, comp129minVal, comp129minI, comp129minJ);
    wire [11:0] comp130minVal;
    wire [5:0] comp130minI, comp130minJ;
    Comparator comp130(SADValues[1030*12 +: 12], 16, 6, SADValues[967*12 +: 12], 15, 7, comp130minVal, comp130minI, comp130minJ);
    wire [11:0] comp131minVal;
    wire [5:0] comp131minI, comp131minJ;
    Comparator comp131(SADValues[904*12 +: 12], 14, 8, SADValues[841*12 +: 12], 13, 9, comp131minVal, comp131minI, comp131minJ);
    wire [11:0] comp132minVal;
    wire [5:0] comp132minI, comp132minJ;
    Comparator comp132(SADValues[778*12 +: 12], 12, 10, SADValues[715*12 +: 12], 11, 11, comp132minVal, comp132minI, comp132minJ);
    wire [11:0] comp133minVal;
    wire [5:0] comp133minI, comp133minJ;
    Comparator comp133(SADValues[652*12 +: 12], 10, 12, SADValues[589*12 +: 12], 9, 13, comp133minVal, comp133minI, comp133minJ);
    wire [11:0] comp134minVal;
    wire [5:0] comp134minI, comp134minJ;
    Comparator comp134(SADValues[526*12 +: 12], 8, 14, SADValues[463*12 +: 12], 7, 15, comp134minVal, comp134minI, comp134minJ);
    wire [11:0] comp135minVal;
    wire [5:0] comp135minI, comp135minJ;
    Comparator comp135(SADValues[400*12 +: 12], 6, 16, SADValues[337*12 +: 12], 5, 17, comp135minVal, comp135minI, comp135minJ);
    wire [11:0] comp136minVal;
    wire [5:0] comp136minI, comp136minJ;
    Comparator comp136(SADValues[274*12 +: 12], 4, 18, SADValues[211*12 +: 12], 3, 19, comp136minVal, comp136minI, comp136minJ);
    wire [11:0] comp137minVal;
    wire [5:0] comp137minI, comp137minJ;
    Comparator comp137(SADValues[148*12 +: 12], 2, 20, SADValues[85*12 +: 12], 1, 21, comp137minVal, comp137minI, comp137minJ);
    wire [11:0] comp138minVal;
    wire [5:0] comp138minI, comp138minJ;
    Comparator comp138(SADValues[22*12 +: 12], 0, 22, SADValues[23*12 +: 12], 0, 23, comp138minVal, comp138minI, comp138minJ);
    wire [11:0] comp139minVal;
    wire [5:0] comp139minI, comp139minJ;
    Comparator comp139(SADValues[86*12 +: 12], 1, 22, SADValues[149*12 +: 12], 2, 21, comp139minVal, comp139minI, comp139minJ);
    wire [11:0] comp140minVal;
    wire [5:0] comp140minI, comp140minJ;
    Comparator comp140(SADValues[212*12 +: 12], 3, 20, SADValues[275*12 +: 12], 4, 19, comp140minVal, comp140minI, comp140minJ);
    wire [11:0] comp141minVal;
    wire [5:0] comp141minI, comp141minJ;
    Comparator comp141(SADValues[338*12 +: 12], 5, 18, SADValues[401*12 +: 12], 6, 17, comp141minVal, comp141minI, comp141minJ);
    wire [11:0] comp142minVal;
    wire [5:0] comp142minI, comp142minJ;
    Comparator comp142(SADValues[464*12 +: 12], 7, 16, SADValues[527*12 +: 12], 8, 15, comp142minVal, comp142minI, comp142minJ);
    wire [11:0] comp143minVal;
    wire [5:0] comp143minI, comp143minJ;
    Comparator comp143(SADValues[590*12 +: 12], 9, 14, SADValues[653*12 +: 12], 10, 13, comp143minVal, comp143minI, comp143minJ);
    wire [11:0] comp144minVal;
    wire [5:0] comp144minI, comp144minJ;
    Comparator comp144(SADValues[716*12 +: 12], 11, 12, SADValues[779*12 +: 12], 12, 11, comp144minVal, comp144minI, comp144minJ);
    wire [11:0] comp145minVal;
    wire [5:0] comp145minI, comp145minJ;
    Comparator comp145(SADValues[842*12 +: 12], 13, 10, SADValues[905*12 +: 12], 14, 9, comp145minVal, comp145minI, comp145minJ);
    wire [11:0] comp146minVal;
    wire [5:0] comp146minI, comp146minJ;
    Comparator comp146(SADValues[968*12 +: 12], 15, 8, SADValues[1031*12 +: 12], 16, 7, comp146minVal, comp146minI, comp146minJ);
    wire [11:0] comp147minVal;
    wire [5:0] comp147minI, comp147minJ;
    Comparator comp147(SADValues[1094*12 +: 12], 17, 6, SADValues[1157*12 +: 12], 18, 5, comp147minVal, comp147minI, comp147minJ);
    wire [11:0] comp148minVal;
    wire [5:0] comp148minI, comp148minJ;
    Comparator comp148(SADValues[1220*12 +: 12], 19, 4, SADValues[1283*12 +: 12], 20, 3, comp148minVal, comp148minI, comp148minJ);
    wire [11:0] comp149minVal;
    wire [5:0] comp149minI, comp149minJ;
    Comparator comp149(SADValues[1346*12 +: 12], 21, 2, SADValues[1409*12 +: 12], 22, 1, comp149minVal, comp149minI, comp149minJ);
    wire [11:0] comp150minVal;
    wire [5:0] comp150minI, comp150minJ;
    Comparator comp150(SADValues[1472*12 +: 12], 23, 0, SADValues[1536*12 +: 12], 24, 0, comp150minVal, comp150minI, comp150minJ);
    wire [11:0] comp151minVal;
    wire [5:0] comp151minI, comp151minJ;
    Comparator comp151(SADValues[1473*12 +: 12], 23, 1, SADValues[1410*12 +: 12], 22, 2, comp151minVal, comp151minI, comp151minJ);
    wire [11:0] comp152minVal;
    wire [5:0] comp152minI, comp152minJ;
    Comparator comp152(SADValues[1347*12 +: 12], 21, 3, SADValues[1284*12 +: 12], 20, 4, comp152minVal, comp152minI, comp152minJ);
    wire [11:0] comp153minVal;
    wire [5:0] comp153minI, comp153minJ;
    Comparator comp153(SADValues[1221*12 +: 12], 19, 5, SADValues[1158*12 +: 12], 18, 6, comp153minVal, comp153minI, comp153minJ);
    wire [11:0] comp154minVal;
    wire [5:0] comp154minI, comp154minJ;
    Comparator comp154(SADValues[1095*12 +: 12], 17, 7, SADValues[1032*12 +: 12], 16, 8, comp154minVal, comp154minI, comp154minJ);
    wire [11:0] comp155minVal;
    wire [5:0] comp155minI, comp155minJ;
    Comparator comp155(SADValues[969*12 +: 12], 15, 9, SADValues[906*12 +: 12], 14, 10, comp155minVal, comp155minI, comp155minJ);
    wire [11:0] comp156minVal;
    wire [5:0] comp156minI, comp156minJ;
    Comparator comp156(SADValues[843*12 +: 12], 13, 11, SADValues[780*12 +: 12], 12, 12, comp156minVal, comp156minI, comp156minJ);
    wire [11:0] comp157minVal;
    wire [5:0] comp157minI, comp157minJ;
    Comparator comp157(SADValues[717*12 +: 12], 11, 13, SADValues[654*12 +: 12], 10, 14, comp157minVal, comp157minI, comp157minJ);
    wire [11:0] comp158minVal;
    wire [5:0] comp158minI, comp158minJ;
    Comparator comp158(SADValues[591*12 +: 12], 9, 15, SADValues[528*12 +: 12], 8, 16, comp158minVal, comp158minI, comp158minJ);
    wire [11:0] comp159minVal;
    wire [5:0] comp159minI, comp159minJ;
    Comparator comp159(SADValues[465*12 +: 12], 7, 17, SADValues[402*12 +: 12], 6, 18, comp159minVal, comp159minI, comp159minJ);
    wire [11:0] comp160minVal;
    wire [5:0] comp160minI, comp160minJ;
    Comparator comp160(SADValues[339*12 +: 12], 5, 19, SADValues[276*12 +: 12], 4, 20, comp160minVal, comp160minI, comp160minJ);
    wire [11:0] comp161minVal;
    wire [5:0] comp161minI, comp161minJ;
    Comparator comp161(SADValues[213*12 +: 12], 3, 21, SADValues[150*12 +: 12], 2, 22, comp161minVal, comp161minI, comp161minJ);
    wire [11:0] comp162minVal;
    wire [5:0] comp162minI, comp162minJ;
    Comparator comp162(SADValues[87*12 +: 12], 1, 23, SADValues[24*12 +: 12], 0, 24, comp162minVal, comp162minI, comp162minJ);
    wire [11:0] comp163minVal;
    wire [5:0] comp163minI, comp163minJ;
    Comparator comp163(SADValues[25*12 +: 12], 0, 25, SADValues[88*12 +: 12], 1, 24, comp163minVal, comp163minI, comp163minJ);
    wire [11:0] comp164minVal;
    wire [5:0] comp164minI, comp164minJ;
    Comparator comp164(SADValues[151*12 +: 12], 2, 23, SADValues[214*12 +: 12], 3, 22, comp164minVal, comp164minI, comp164minJ);
    wire [11:0] comp165minVal;
    wire [5:0] comp165minI, comp165minJ;
    Comparator comp165(SADValues[277*12 +: 12], 4, 21, SADValues[340*12 +: 12], 5, 20, comp165minVal, comp165minI, comp165minJ);
    wire [11:0] comp166minVal;
    wire [5:0] comp166minI, comp166minJ;
    Comparator comp166(SADValues[403*12 +: 12], 6, 19, SADValues[466*12 +: 12], 7, 18, comp166minVal, comp166minI, comp166minJ);
    wire [11:0] comp167minVal;
    wire [5:0] comp167minI, comp167minJ;
    Comparator comp167(SADValues[529*12 +: 12], 8, 17, SADValues[592*12 +: 12], 9, 16, comp167minVal, comp167minI, comp167minJ);
    wire [11:0] comp168minVal;
    wire [5:0] comp168minI, comp168minJ;
    Comparator comp168(SADValues[655*12 +: 12], 10, 15, SADValues[718*12 +: 12], 11, 14, comp168minVal, comp168minI, comp168minJ);
    wire [11:0] comp169minVal;
    wire [5:0] comp169minI, comp169minJ;
    Comparator comp169(SADValues[781*12 +: 12], 12, 13, SADValues[844*12 +: 12], 13, 12, comp169minVal, comp169minI, comp169minJ);
    wire [11:0] comp170minVal;
    wire [5:0] comp170minI, comp170minJ;
    Comparator comp170(SADValues[907*12 +: 12], 14, 11, SADValues[970*12 +: 12], 15, 10, comp170minVal, comp170minI, comp170minJ);
    wire [11:0] comp171minVal;
    wire [5:0] comp171minI, comp171minJ;
    Comparator comp171(SADValues[1033*12 +: 12], 16, 9, SADValues[1096*12 +: 12], 17, 8, comp171minVal, comp171minI, comp171minJ);
    wire [11:0] comp172minVal;
    wire [5:0] comp172minI, comp172minJ;
    Comparator comp172(SADValues[1159*12 +: 12], 18, 7, SADValues[1222*12 +: 12], 19, 6, comp172minVal, comp172minI, comp172minJ);
    wire [11:0] comp173minVal;
    wire [5:0] comp173minI, comp173minJ;
    Comparator comp173(SADValues[1285*12 +: 12], 20, 5, SADValues[1348*12 +: 12], 21, 4, comp173minVal, comp173minI, comp173minJ);
    wire [11:0] comp174minVal;
    wire [5:0] comp174minI, comp174minJ;
    Comparator comp174(SADValues[1411*12 +: 12], 22, 3, SADValues[1474*12 +: 12], 23, 2, comp174minVal, comp174minI, comp174minJ);
    wire [11:0] comp175minVal;
    wire [5:0] comp175minI, comp175minJ;
    Comparator comp175(SADValues[1537*12 +: 12], 24, 1, SADValues[1600*12 +: 12], 25, 0, comp175minVal, comp175minI, comp175minJ);
    wire [11:0] comp176minVal;
    wire [5:0] comp176minI, comp176minJ;
    Comparator comp176(SADValues[1664*12 +: 12], 26, 0, SADValues[1601*12 +: 12], 25, 1, comp176minVal, comp176minI, comp176minJ);
    wire [11:0] comp177minVal;
    wire [5:0] comp177minI, comp177minJ;
    Comparator comp177(SADValues[1538*12 +: 12], 24, 2, SADValues[1475*12 +: 12], 23, 3, comp177minVal, comp177minI, comp177minJ);
    wire [11:0] comp178minVal;
    wire [5:0] comp178minI, comp178minJ;
    Comparator comp178(SADValues[1412*12 +: 12], 22, 4, SADValues[1349*12 +: 12], 21, 5, comp178minVal, comp178minI, comp178minJ);
    wire [11:0] comp179minVal;
    wire [5:0] comp179minI, comp179minJ;
    Comparator comp179(SADValues[1286*12 +: 12], 20, 6, SADValues[1223*12 +: 12], 19, 7, comp179minVal, comp179minI, comp179minJ);
    wire [11:0] comp180minVal;
    wire [5:0] comp180minI, comp180minJ;
    Comparator comp180(SADValues[1160*12 +: 12], 18, 8, SADValues[1097*12 +: 12], 17, 9, comp180minVal, comp180minI, comp180minJ);
    wire [11:0] comp181minVal;
    wire [5:0] comp181minI, comp181minJ;
    Comparator comp181(SADValues[1034*12 +: 12], 16, 10, SADValues[971*12 +: 12], 15, 11, comp181minVal, comp181minI, comp181minJ);
    wire [11:0] comp182minVal;
    wire [5:0] comp182minI, comp182minJ;
    Comparator comp182(SADValues[908*12 +: 12], 14, 12, SADValues[845*12 +: 12], 13, 13, comp182minVal, comp182minI, comp182minJ);
    wire [11:0] comp183minVal;
    wire [5:0] comp183minI, comp183minJ;
    Comparator comp183(SADValues[782*12 +: 12], 12, 14, SADValues[719*12 +: 12], 11, 15, comp183minVal, comp183minI, comp183minJ);
    wire [11:0] comp184minVal;
    wire [5:0] comp184minI, comp184minJ;
    Comparator comp184(SADValues[656*12 +: 12], 10, 16, SADValues[593*12 +: 12], 9, 17, comp184minVal, comp184minI, comp184minJ);
    wire [11:0] comp185minVal;
    wire [5:0] comp185minI, comp185minJ;
    Comparator comp185(SADValues[530*12 +: 12], 8, 18, SADValues[467*12 +: 12], 7, 19, comp185minVal, comp185minI, comp185minJ);
    wire [11:0] comp186minVal;
    wire [5:0] comp186minI, comp186minJ;
    Comparator comp186(SADValues[404*12 +: 12], 6, 20, SADValues[341*12 +: 12], 5, 21, comp186minVal, comp186minI, comp186minJ);
    wire [11:0] comp187minVal;
    wire [5:0] comp187minI, comp187minJ;
    Comparator comp187(SADValues[278*12 +: 12], 4, 22, SADValues[215*12 +: 12], 3, 23, comp187minVal, comp187minI, comp187minJ);
    wire [11:0] comp188minVal;
    wire [5:0] comp188minI, comp188minJ;
    Comparator comp188(SADValues[152*12 +: 12], 2, 24, SADValues[89*12 +: 12], 1, 25, comp188minVal, comp188minI, comp188minJ);
    wire [11:0] comp189minVal;
    wire [5:0] comp189minI, comp189minJ;
    Comparator comp189(SADValues[26*12 +: 12], 0, 26, SADValues[27*12 +: 12], 0, 27, comp189minVal, comp189minI, comp189minJ);
    wire [11:0] comp190minVal;
    wire [5:0] comp190minI, comp190minJ;
    Comparator comp190(SADValues[90*12 +: 12], 1, 26, SADValues[153*12 +: 12], 2, 25, comp190minVal, comp190minI, comp190minJ);
    wire [11:0] comp191minVal;
    wire [5:0] comp191minI, comp191minJ;
    Comparator comp191(SADValues[216*12 +: 12], 3, 24, SADValues[279*12 +: 12], 4, 23, comp191minVal, comp191minI, comp191minJ);
    wire [11:0] comp192minVal;
    wire [5:0] comp192minI, comp192minJ;
    Comparator comp192(SADValues[342*12 +: 12], 5, 22, SADValues[405*12 +: 12], 6, 21, comp192minVal, comp192minI, comp192minJ);
    wire [11:0] comp193minVal;
    wire [5:0] comp193minI, comp193minJ;
    Comparator comp193(SADValues[468*12 +: 12], 7, 20, SADValues[531*12 +: 12], 8, 19, comp193minVal, comp193minI, comp193minJ);
    wire [11:0] comp194minVal;
    wire [5:0] comp194minI, comp194minJ;
    Comparator comp194(SADValues[594*12 +: 12], 9, 18, SADValues[657*12 +: 12], 10, 17, comp194minVal, comp194minI, comp194minJ);
    wire [11:0] comp195minVal;
    wire [5:0] comp195minI, comp195minJ;
    Comparator comp195(SADValues[720*12 +: 12], 11, 16, SADValues[783*12 +: 12], 12, 15, comp195minVal, comp195minI, comp195minJ);
    wire [11:0] comp196minVal;
    wire [5:0] comp196minI, comp196minJ;
    Comparator comp196(SADValues[846*12 +: 12], 13, 14, SADValues[909*12 +: 12], 14, 13, comp196minVal, comp196minI, comp196minJ);
    wire [11:0] comp197minVal;
    wire [5:0] comp197minI, comp197minJ;
    Comparator comp197(SADValues[972*12 +: 12], 15, 12, SADValues[1035*12 +: 12], 16, 11, comp197minVal, comp197minI, comp197minJ);
    wire [11:0] comp198minVal;
    wire [5:0] comp198minI, comp198minJ;
    Comparator comp198(SADValues[1098*12 +: 12], 17, 10, SADValues[1161*12 +: 12], 18, 9, comp198minVal, comp198minI, comp198minJ);
    wire [11:0] comp199minVal;
    wire [5:0] comp199minI, comp199minJ;
    Comparator comp199(SADValues[1224*12 +: 12], 19, 8, SADValues[1287*12 +: 12], 20, 7, comp199minVal, comp199minI, comp199minJ);
    wire [11:0] comp200minVal;
    wire [5:0] comp200minI, comp200minJ;
    Comparator comp200(SADValues[1350*12 +: 12], 21, 6, SADValues[1413*12 +: 12], 22, 5, comp200minVal, comp200minI, comp200minJ);
    wire [11:0] comp201minVal;
    wire [5:0] comp201minI, comp201minJ;
    Comparator comp201(SADValues[1476*12 +: 12], 23, 4, SADValues[1539*12 +: 12], 24, 3, comp201minVal, comp201minI, comp201minJ);
    wire [11:0] comp202minVal;
    wire [5:0] comp202minI, comp202minJ;
    Comparator comp202(SADValues[1602*12 +: 12], 25, 2, SADValues[1665*12 +: 12], 26, 1, comp202minVal, comp202minI, comp202minJ);
    wire [11:0] comp203minVal;
    wire [5:0] comp203minI, comp203minJ;
    Comparator comp203(SADValues[1728*12 +: 12], 27, 0, SADValues[1792*12 +: 12], 28, 0, comp203minVal, comp203minI, comp203minJ);
    wire [11:0] comp204minVal;
    wire [5:0] comp204minI, comp204minJ;
    Comparator comp204(SADValues[1729*12 +: 12], 27, 1, SADValues[1666*12 +: 12], 26, 2, comp204minVal, comp204minI, comp204minJ);
    wire [11:0] comp205minVal;
    wire [5:0] comp205minI, comp205minJ;
    Comparator comp205(SADValues[1603*12 +: 12], 25, 3, SADValues[1540*12 +: 12], 24, 4, comp205minVal, comp205minI, comp205minJ);
    wire [11:0] comp206minVal;
    wire [5:0] comp206minI, comp206minJ;
    Comparator comp206(SADValues[1477*12 +: 12], 23, 5, SADValues[1414*12 +: 12], 22, 6, comp206minVal, comp206minI, comp206minJ);
    wire [11:0] comp207minVal;
    wire [5:0] comp207minI, comp207minJ;
    Comparator comp207(SADValues[1351*12 +: 12], 21, 7, SADValues[1288*12 +: 12], 20, 8, comp207minVal, comp207minI, comp207minJ);
    wire [11:0] comp208minVal;
    wire [5:0] comp208minI, comp208minJ;
    Comparator comp208(SADValues[1225*12 +: 12], 19, 9, SADValues[1162*12 +: 12], 18, 10, comp208minVal, comp208minI, comp208minJ);
    wire [11:0] comp209minVal;
    wire [5:0] comp209minI, comp209minJ;
    Comparator comp209(SADValues[1099*12 +: 12], 17, 11, SADValues[1036*12 +: 12], 16, 12, comp209minVal, comp209minI, comp209minJ);
    wire [11:0] comp210minVal;
    wire [5:0] comp210minI, comp210minJ;
    Comparator comp210(SADValues[973*12 +: 12], 15, 13, SADValues[910*12 +: 12], 14, 14, comp210minVal, comp210minI, comp210minJ);
    wire [11:0] comp211minVal;
    wire [5:0] comp211minI, comp211minJ;
    Comparator comp211(SADValues[847*12 +: 12], 13, 15, SADValues[784*12 +: 12], 12, 16, comp211minVal, comp211minI, comp211minJ);
    wire [11:0] comp212minVal;
    wire [5:0] comp212minI, comp212minJ;
    Comparator comp212(SADValues[721*12 +: 12], 11, 17, SADValues[658*12 +: 12], 10, 18, comp212minVal, comp212minI, comp212minJ);
    wire [11:0] comp213minVal;
    wire [5:0] comp213minI, comp213minJ;
    Comparator comp213(SADValues[595*12 +: 12], 9, 19, SADValues[532*12 +: 12], 8, 20, comp213minVal, comp213minI, comp213minJ);
    wire [11:0] comp214minVal;
    wire [5:0] comp214minI, comp214minJ;
    Comparator comp214(SADValues[469*12 +: 12], 7, 21, SADValues[406*12 +: 12], 6, 22, comp214minVal, comp214minI, comp214minJ);
    wire [11:0] comp215minVal;
    wire [5:0] comp215minI, comp215minJ;
    Comparator comp215(SADValues[343*12 +: 12], 5, 23, SADValues[280*12 +: 12], 4, 24, comp215minVal, comp215minI, comp215minJ);
    wire [11:0] comp216minVal;
    wire [5:0] comp216minI, comp216minJ;
    Comparator comp216(SADValues[217*12 +: 12], 3, 25, SADValues[154*12 +: 12], 2, 26, comp216minVal, comp216minI, comp216minJ);
    wire [11:0] comp217minVal;
    wire [5:0] comp217minI, comp217minJ;
    Comparator comp217(SADValues[91*12 +: 12], 1, 27, SADValues[28*12 +: 12], 0, 28, comp217minVal, comp217minI, comp217minJ);
    wire [11:0] comp218minVal;
    wire [5:0] comp218minI, comp218minJ;
    Comparator comp218(SADValues[29*12 +: 12], 0, 29, SADValues[92*12 +: 12], 1, 28, comp218minVal, comp218minI, comp218minJ);
    wire [11:0] comp219minVal;
    wire [5:0] comp219minI, comp219minJ;
    Comparator comp219(SADValues[155*12 +: 12], 2, 27, SADValues[218*12 +: 12], 3, 26, comp219minVal, comp219minI, comp219minJ);
    wire [11:0] comp220minVal;
    wire [5:0] comp220minI, comp220minJ;
    Comparator comp220(SADValues[281*12 +: 12], 4, 25, SADValues[344*12 +: 12], 5, 24, comp220minVal, comp220minI, comp220minJ);
    wire [11:0] comp221minVal;
    wire [5:0] comp221minI, comp221minJ;
    Comparator comp221(SADValues[407*12 +: 12], 6, 23, SADValues[470*12 +: 12], 7, 22, comp221minVal, comp221minI, comp221minJ);
    wire [11:0] comp222minVal;
    wire [5:0] comp222minI, comp222minJ;
    Comparator comp222(SADValues[533*12 +: 12], 8, 21, SADValues[596*12 +: 12], 9, 20, comp222minVal, comp222minI, comp222minJ);
    wire [11:0] comp223minVal;
    wire [5:0] comp223minI, comp223minJ;
    Comparator comp223(SADValues[659*12 +: 12], 10, 19, SADValues[722*12 +: 12], 11, 18, comp223minVal, comp223minI, comp223minJ);
    wire [11:0] comp224minVal;
    wire [5:0] comp224minI, comp224minJ;
    Comparator comp224(SADValues[785*12 +: 12], 12, 17, SADValues[848*12 +: 12], 13, 16, comp224minVal, comp224minI, comp224minJ);
    wire [11:0] comp225minVal;
    wire [5:0] comp225minI, comp225minJ;
    Comparator comp225(SADValues[911*12 +: 12], 14, 15, SADValues[974*12 +: 12], 15, 14, comp225minVal, comp225minI, comp225minJ);
    wire [11:0] comp226minVal;
    wire [5:0] comp226minI, comp226minJ;
    Comparator comp226(SADValues[1037*12 +: 12], 16, 13, SADValues[1100*12 +: 12], 17, 12, comp226minVal, comp226minI, comp226minJ);
    wire [11:0] comp227minVal;
    wire [5:0] comp227minI, comp227minJ;
    Comparator comp227(SADValues[1163*12 +: 12], 18, 11, SADValues[1226*12 +: 12], 19, 10, comp227minVal, comp227minI, comp227minJ);
    wire [11:0] comp228minVal;
    wire [5:0] comp228minI, comp228minJ;
    Comparator comp228(SADValues[1289*12 +: 12], 20, 9, SADValues[1352*12 +: 12], 21, 8, comp228minVal, comp228minI, comp228minJ);
    wire [11:0] comp229minVal;
    wire [5:0] comp229minI, comp229minJ;
    Comparator comp229(SADValues[1415*12 +: 12], 22, 7, SADValues[1478*12 +: 12], 23, 6, comp229minVal, comp229minI, comp229minJ);
    wire [11:0] comp230minVal;
    wire [5:0] comp230minI, comp230minJ;
    Comparator comp230(SADValues[1541*12 +: 12], 24, 5, SADValues[1604*12 +: 12], 25, 4, comp230minVal, comp230minI, comp230minJ);
    wire [11:0] comp231minVal;
    wire [5:0] comp231minI, comp231minJ;
    Comparator comp231(SADValues[1667*12 +: 12], 26, 3, SADValues[1730*12 +: 12], 27, 2, comp231minVal, comp231minI, comp231minJ);
    wire [11:0] comp232minVal;
    wire [5:0] comp232minI, comp232minJ;
    Comparator comp232(SADValues[1793*12 +: 12], 28, 1, SADValues[1856*12 +: 12], 29, 0, comp232minVal, comp232minI, comp232minJ);
    wire [11:0] comp233minVal;
    wire [5:0] comp233minI, comp233minJ;
    Comparator comp233(SADValues[1920*12 +: 12], 30, 0, SADValues[1857*12 +: 12], 29, 1, comp233minVal, comp233minI, comp233minJ);
    wire [11:0] comp234minVal;
    wire [5:0] comp234minI, comp234minJ;
    Comparator comp234(SADValues[1794*12 +: 12], 28, 2, SADValues[1731*12 +: 12], 27, 3, comp234minVal, comp234minI, comp234minJ);
    wire [11:0] comp235minVal;
    wire [5:0] comp235minI, comp235minJ;
    Comparator comp235(SADValues[1668*12 +: 12], 26, 4, SADValues[1605*12 +: 12], 25, 5, comp235minVal, comp235minI, comp235minJ);
    wire [11:0] comp236minVal;
    wire [5:0] comp236minI, comp236minJ;
    Comparator comp236(SADValues[1542*12 +: 12], 24, 6, SADValues[1479*12 +: 12], 23, 7, comp236minVal, comp236minI, comp236minJ);
    wire [11:0] comp237minVal;
    wire [5:0] comp237minI, comp237minJ;
    Comparator comp237(SADValues[1416*12 +: 12], 22, 8, SADValues[1353*12 +: 12], 21, 9, comp237minVal, comp237minI, comp237minJ);
    wire [11:0] comp238minVal;
    wire [5:0] comp238minI, comp238minJ;
    Comparator comp238(SADValues[1290*12 +: 12], 20, 10, SADValues[1227*12 +: 12], 19, 11, comp238minVal, comp238minI, comp238minJ);
    wire [11:0] comp239minVal;
    wire [5:0] comp239minI, comp239minJ;
    Comparator comp239(SADValues[1164*12 +: 12], 18, 12, SADValues[1101*12 +: 12], 17, 13, comp239minVal, comp239minI, comp239minJ);
    wire [11:0] comp240minVal;
    wire [5:0] comp240minI, comp240minJ;
    Comparator comp240(SADValues[1038*12 +: 12], 16, 14, SADValues[975*12 +: 12], 15, 15, comp240minVal, comp240minI, comp240minJ);
    wire [11:0] comp241minVal;
    wire [5:0] comp241minI, comp241minJ;
    Comparator comp241(SADValues[912*12 +: 12], 14, 16, SADValues[849*12 +: 12], 13, 17, comp241minVal, comp241minI, comp241minJ);
    wire [11:0] comp242minVal;
    wire [5:0] comp242minI, comp242minJ;
    Comparator comp242(SADValues[786*12 +: 12], 12, 18, SADValues[723*12 +: 12], 11, 19, comp242minVal, comp242minI, comp242minJ);
    wire [11:0] comp243minVal;
    wire [5:0] comp243minI, comp243minJ;
    Comparator comp243(SADValues[660*12 +: 12], 10, 20, SADValues[597*12 +: 12], 9, 21, comp243minVal, comp243minI, comp243minJ);
    wire [11:0] comp244minVal;
    wire [5:0] comp244minI, comp244minJ;
    Comparator comp244(SADValues[534*12 +: 12], 8, 22, SADValues[471*12 +: 12], 7, 23, comp244minVal, comp244minI, comp244minJ);
    wire [11:0] comp245minVal;
    wire [5:0] comp245minI, comp245minJ;
    Comparator comp245(SADValues[408*12 +: 12], 6, 24, SADValues[345*12 +: 12], 5, 25, comp245minVal, comp245minI, comp245minJ);
    wire [11:0] comp246minVal;
    wire [5:0] comp246minI, comp246minJ;
    Comparator comp246(SADValues[282*12 +: 12], 4, 26, SADValues[219*12 +: 12], 3, 27, comp246minVal, comp246minI, comp246minJ);
    wire [11:0] comp247minVal;
    wire [5:0] comp247minI, comp247minJ;
    Comparator comp247(SADValues[156*12 +: 12], 2, 28, SADValues[93*12 +: 12], 1, 29, comp247minVal, comp247minI, comp247minJ);
    wire [11:0] comp248minVal;
    wire [5:0] comp248minI, comp248minJ;
    Comparator comp248(SADValues[30*12 +: 12], 0, 30, SADValues[31*12 +: 12], 0, 31, comp248minVal, comp248minI, comp248minJ);
    wire [11:0] comp249minVal;
    wire [5:0] comp249minI, comp249minJ;
    Comparator comp249(SADValues[94*12 +: 12], 1, 30, SADValues[157*12 +: 12], 2, 29, comp249minVal, comp249minI, comp249minJ);
    wire [11:0] comp250minVal;
    wire [5:0] comp250minI, comp250minJ;
    Comparator comp250(SADValues[220*12 +: 12], 3, 28, SADValues[283*12 +: 12], 4, 27, comp250minVal, comp250minI, comp250minJ);
    wire [11:0] comp251minVal;
    wire [5:0] comp251minI, comp251minJ;
    Comparator comp251(SADValues[346*12 +: 12], 5, 26, SADValues[409*12 +: 12], 6, 25, comp251minVal, comp251minI, comp251minJ);
    wire [11:0] comp252minVal;
    wire [5:0] comp252minI, comp252minJ;
    Comparator comp252(SADValues[472*12 +: 12], 7, 24, SADValues[535*12 +: 12], 8, 23, comp252minVal, comp252minI, comp252minJ);
    wire [11:0] comp253minVal;
    wire [5:0] comp253minI, comp253minJ;
    Comparator comp253(SADValues[598*12 +: 12], 9, 22, SADValues[661*12 +: 12], 10, 21, comp253minVal, comp253minI, comp253minJ);
    wire [11:0] comp254minVal;
    wire [5:0] comp254minI, comp254minJ;
    Comparator comp254(SADValues[724*12 +: 12], 11, 20, SADValues[787*12 +: 12], 12, 19, comp254minVal, comp254minI, comp254minJ);
    wire [11:0] comp255minVal;
    wire [5:0] comp255minI, comp255minJ;
    Comparator comp255(SADValues[850*12 +: 12], 13, 18, SADValues[913*12 +: 12], 14, 17, comp255minVal, comp255minI, comp255minJ);
    wire [11:0] comp256minVal;
    wire [5:0] comp256minI, comp256minJ;
    Comparator comp256(SADValues[976*12 +: 12], 15, 16, SADValues[1039*12 +: 12], 16, 15, comp256minVal, comp256minI, comp256minJ);
    wire [11:0] comp257minVal;
    wire [5:0] comp257minI, comp257minJ;
    Comparator comp257(SADValues[1102*12 +: 12], 17, 14, SADValues[1165*12 +: 12], 18, 13, comp257minVal, comp257minI, comp257minJ);
    wire [11:0] comp258minVal;
    wire [5:0] comp258minI, comp258minJ;
    Comparator comp258(SADValues[1228*12 +: 12], 19, 12, SADValues[1291*12 +: 12], 20, 11, comp258minVal, comp258minI, comp258minJ);
    wire [11:0] comp259minVal;
    wire [5:0] comp259minI, comp259minJ;
    Comparator comp259(SADValues[1354*12 +: 12], 21, 10, SADValues[1417*12 +: 12], 22, 9, comp259minVal, comp259minI, comp259minJ);
    wire [11:0] comp260minVal;
    wire [5:0] comp260minI, comp260minJ;
    Comparator comp260(SADValues[1480*12 +: 12], 23, 8, SADValues[1543*12 +: 12], 24, 7, comp260minVal, comp260minI, comp260minJ);
    wire [11:0] comp261minVal;
    wire [5:0] comp261minI, comp261minJ;
    Comparator comp261(SADValues[1606*12 +: 12], 25, 6, SADValues[1669*12 +: 12], 26, 5, comp261minVal, comp261minI, comp261minJ);
    wire [11:0] comp262minVal;
    wire [5:0] comp262minI, comp262minJ;
    Comparator comp262(SADValues[1732*12 +: 12], 27, 4, SADValues[1795*12 +: 12], 28, 3, comp262minVal, comp262minI, comp262minJ);
    wire [11:0] comp263minVal;
    wire [5:0] comp263minI, comp263minJ;
    Comparator comp263(SADValues[1858*12 +: 12], 29, 2, SADValues[1921*12 +: 12], 30, 1, comp263minVal, comp263minI, comp263minJ);
    wire [11:0] comp264minVal;
    wire [5:0] comp264minI, comp264minJ;
    Comparator comp264(SADValues[1984*12 +: 12], 31, 0, SADValues[2048*12 +: 12], 32, 0, comp264minVal, comp264minI, comp264minJ);
    wire [11:0] comp265minVal;
    wire [5:0] comp265minI, comp265minJ;
    Comparator comp265(SADValues[1985*12 +: 12], 31, 1, SADValues[1922*12 +: 12], 30, 2, comp265minVal, comp265minI, comp265minJ);
    wire [11:0] comp266minVal;
    wire [5:0] comp266minI, comp266minJ;
    Comparator comp266(SADValues[1859*12 +: 12], 29, 3, SADValues[1796*12 +: 12], 28, 4, comp266minVal, comp266minI, comp266minJ);
    wire [11:0] comp267minVal;
    wire [5:0] comp267minI, comp267minJ;
    Comparator comp267(SADValues[1733*12 +: 12], 27, 5, SADValues[1670*12 +: 12], 26, 6, comp267minVal, comp267minI, comp267minJ);
    wire [11:0] comp268minVal;
    wire [5:0] comp268minI, comp268minJ;
    Comparator comp268(SADValues[1607*12 +: 12], 25, 7, SADValues[1544*12 +: 12], 24, 8, comp268minVal, comp268minI, comp268minJ);
    wire [11:0] comp269minVal;
    wire [5:0] comp269minI, comp269minJ;
    Comparator comp269(SADValues[1481*12 +: 12], 23, 9, SADValues[1418*12 +: 12], 22, 10, comp269minVal, comp269minI, comp269minJ);
    wire [11:0] comp270minVal;
    wire [5:0] comp270minI, comp270minJ;
    Comparator comp270(SADValues[1355*12 +: 12], 21, 11, SADValues[1292*12 +: 12], 20, 12, comp270minVal, comp270minI, comp270minJ);
    wire [11:0] comp271minVal;
    wire [5:0] comp271minI, comp271minJ;
    Comparator comp271(SADValues[1229*12 +: 12], 19, 13, SADValues[1166*12 +: 12], 18, 14, comp271minVal, comp271minI, comp271minJ);
    wire [11:0] comp272minVal;
    wire [5:0] comp272minI, comp272minJ;
    Comparator comp272(SADValues[1103*12 +: 12], 17, 15, SADValues[1040*12 +: 12], 16, 16, comp272minVal, comp272minI, comp272minJ);
    wire [11:0] comp273minVal;
    wire [5:0] comp273minI, comp273minJ;
    Comparator comp273(SADValues[977*12 +: 12], 15, 17, SADValues[914*12 +: 12], 14, 18, comp273minVal, comp273minI, comp273minJ);
    wire [11:0] comp274minVal;
    wire [5:0] comp274minI, comp274minJ;
    Comparator comp274(SADValues[851*12 +: 12], 13, 19, SADValues[788*12 +: 12], 12, 20, comp274minVal, comp274minI, comp274minJ);
    wire [11:0] comp275minVal;
    wire [5:0] comp275minI, comp275minJ;
    Comparator comp275(SADValues[725*12 +: 12], 11, 21, SADValues[662*12 +: 12], 10, 22, comp275minVal, comp275minI, comp275minJ);
    wire [11:0] comp276minVal;
    wire [5:0] comp276minI, comp276minJ;
    Comparator comp276(SADValues[599*12 +: 12], 9, 23, SADValues[536*12 +: 12], 8, 24, comp276minVal, comp276minI, comp276minJ);
    wire [11:0] comp277minVal;
    wire [5:0] comp277minI, comp277minJ;
    Comparator comp277(SADValues[473*12 +: 12], 7, 25, SADValues[410*12 +: 12], 6, 26, comp277minVal, comp277minI, comp277minJ);
    wire [11:0] comp278minVal;
    wire [5:0] comp278minI, comp278minJ;
    Comparator comp278(SADValues[347*12 +: 12], 5, 27, SADValues[284*12 +: 12], 4, 28, comp278minVal, comp278minI, comp278minJ);
    wire [11:0] comp279minVal;
    wire [5:0] comp279minI, comp279minJ;
    Comparator comp279(SADValues[221*12 +: 12], 3, 29, SADValues[158*12 +: 12], 2, 30, comp279minVal, comp279minI, comp279minJ);
    wire [11:0] comp280minVal;
    wire [5:0] comp280minI, comp280minJ;
    Comparator comp280(SADValues[95*12 +: 12], 1, 31, SADValues[32*12 +: 12], 0, 32, comp280minVal, comp280minI, comp280minJ);
    wire [11:0] comp281minVal;
    wire [5:0] comp281minI, comp281minJ;
    Comparator comp281(SADValues[33*12 +: 12], 0, 33, SADValues[96*12 +: 12], 1, 32, comp281minVal, comp281minI, comp281minJ);
    wire [11:0] comp282minVal;
    wire [5:0] comp282minI, comp282minJ;
    Comparator comp282(SADValues[159*12 +: 12], 2, 31, SADValues[222*12 +: 12], 3, 30, comp282minVal, comp282minI, comp282minJ);
    wire [11:0] comp283minVal;
    wire [5:0] comp283minI, comp283minJ;
    Comparator comp283(SADValues[285*12 +: 12], 4, 29, SADValues[348*12 +: 12], 5, 28, comp283minVal, comp283minI, comp283minJ);
    wire [11:0] comp284minVal;
    wire [5:0] comp284minI, comp284minJ;
    Comparator comp284(SADValues[411*12 +: 12], 6, 27, SADValues[474*12 +: 12], 7, 26, comp284minVal, comp284minI, comp284minJ);
    wire [11:0] comp285minVal;
    wire [5:0] comp285minI, comp285minJ;
    Comparator comp285(SADValues[537*12 +: 12], 8, 25, SADValues[600*12 +: 12], 9, 24, comp285minVal, comp285minI, comp285minJ);
    wire [11:0] comp286minVal;
    wire [5:0] comp286minI, comp286minJ;
    Comparator comp286(SADValues[663*12 +: 12], 10, 23, SADValues[726*12 +: 12], 11, 22, comp286minVal, comp286minI, comp286minJ);
    wire [11:0] comp287minVal;
    wire [5:0] comp287minI, comp287minJ;
    Comparator comp287(SADValues[789*12 +: 12], 12, 21, SADValues[852*12 +: 12], 13, 20, comp287minVal, comp287minI, comp287minJ);
    wire [11:0] comp288minVal;
    wire [5:0] comp288minI, comp288minJ;
    Comparator comp288(SADValues[915*12 +: 12], 14, 19, SADValues[978*12 +: 12], 15, 18, comp288minVal, comp288minI, comp288minJ);
    wire [11:0] comp289minVal;
    wire [5:0] comp289minI, comp289minJ;
    Comparator comp289(SADValues[1041*12 +: 12], 16, 17, SADValues[1104*12 +: 12], 17, 16, comp289minVal, comp289minI, comp289minJ);
    wire [11:0] comp290minVal;
    wire [5:0] comp290minI, comp290minJ;
    Comparator comp290(SADValues[1167*12 +: 12], 18, 15, SADValues[1230*12 +: 12], 19, 14, comp290minVal, comp290minI, comp290minJ);
    wire [11:0] comp291minVal;
    wire [5:0] comp291minI, comp291minJ;
    Comparator comp291(SADValues[1293*12 +: 12], 20, 13, SADValues[1356*12 +: 12], 21, 12, comp291minVal, comp291minI, comp291minJ);
    wire [11:0] comp292minVal;
    wire [5:0] comp292minI, comp292minJ;
    Comparator comp292(SADValues[1419*12 +: 12], 22, 11, SADValues[1482*12 +: 12], 23, 10, comp292minVal, comp292minI, comp292minJ);
    wire [11:0] comp293minVal;
    wire [5:0] comp293minI, comp293minJ;
    Comparator comp293(SADValues[1545*12 +: 12], 24, 9, SADValues[1608*12 +: 12], 25, 8, comp293minVal, comp293minI, comp293minJ);
    wire [11:0] comp294minVal;
    wire [5:0] comp294minI, comp294minJ;
    Comparator comp294(SADValues[1671*12 +: 12], 26, 7, SADValues[1734*12 +: 12], 27, 6, comp294minVal, comp294minI, comp294minJ);
    wire [11:0] comp295minVal;
    wire [5:0] comp295minI, comp295minJ;
    Comparator comp295(SADValues[1797*12 +: 12], 28, 5, SADValues[1860*12 +: 12], 29, 4, comp295minVal, comp295minI, comp295minJ);
    wire [11:0] comp296minVal;
    wire [5:0] comp296minI, comp296minJ;
    Comparator comp296(SADValues[1923*12 +: 12], 30, 3, SADValues[1986*12 +: 12], 31, 2, comp296minVal, comp296minI, comp296minJ);
    wire [11:0] comp297minVal;
    wire [5:0] comp297minI, comp297minJ;
    Comparator comp297(SADValues[2049*12 +: 12], 32, 1, SADValues[2112*12 +: 12], 33, 0, comp297minVal, comp297minI, comp297minJ);
    wire [11:0] comp298minVal;
    wire [5:0] comp298minI, comp298minJ;
    Comparator comp298(SADValues[2176*12 +: 12], 34, 0, SADValues[2113*12 +: 12], 33, 1, comp298minVal, comp298minI, comp298minJ);
    wire [11:0] comp299minVal;
    wire [5:0] comp299minI, comp299minJ;
    Comparator comp299(SADValues[2050*12 +: 12], 32, 2, SADValues[1987*12 +: 12], 31, 3, comp299minVal, comp299minI, comp299minJ);
    wire [11:0] comp300minVal;
    wire [5:0] comp300minI, comp300minJ;
    Comparator comp300(SADValues[1924*12 +: 12], 30, 4, SADValues[1861*12 +: 12], 29, 5, comp300minVal, comp300minI, comp300minJ);
    wire [11:0] comp301minVal;
    wire [5:0] comp301minI, comp301minJ;
    Comparator comp301(SADValues[1798*12 +: 12], 28, 6, SADValues[1735*12 +: 12], 27, 7, comp301minVal, comp301minI, comp301minJ);
    wire [11:0] comp302minVal;
    wire [5:0] comp302minI, comp302minJ;
    Comparator comp302(SADValues[1672*12 +: 12], 26, 8, SADValues[1609*12 +: 12], 25, 9, comp302minVal, comp302minI, comp302minJ);
    wire [11:0] comp303minVal;
    wire [5:0] comp303minI, comp303minJ;
    Comparator comp303(SADValues[1546*12 +: 12], 24, 10, SADValues[1483*12 +: 12], 23, 11, comp303minVal, comp303minI, comp303minJ);
    wire [11:0] comp304minVal;
    wire [5:0] comp304minI, comp304minJ;
    Comparator comp304(SADValues[1420*12 +: 12], 22, 12, SADValues[1357*12 +: 12], 21, 13, comp304minVal, comp304minI, comp304minJ);
    wire [11:0] comp305minVal;
    wire [5:0] comp305minI, comp305minJ;
    Comparator comp305(SADValues[1294*12 +: 12], 20, 14, SADValues[1231*12 +: 12], 19, 15, comp305minVal, comp305minI, comp305minJ);
    wire [11:0] comp306minVal;
    wire [5:0] comp306minI, comp306minJ;
    Comparator comp306(SADValues[1168*12 +: 12], 18, 16, SADValues[1105*12 +: 12], 17, 17, comp306minVal, comp306minI, comp306minJ);
    wire [11:0] comp307minVal;
    wire [5:0] comp307minI, comp307minJ;
    Comparator comp307(SADValues[1042*12 +: 12], 16, 18, SADValues[979*12 +: 12], 15, 19, comp307minVal, comp307minI, comp307minJ);
    wire [11:0] comp308minVal;
    wire [5:0] comp308minI, comp308minJ;
    Comparator comp308(SADValues[916*12 +: 12], 14, 20, SADValues[853*12 +: 12], 13, 21, comp308minVal, comp308minI, comp308minJ);
    wire [11:0] comp309minVal;
    wire [5:0] comp309minI, comp309minJ;
    Comparator comp309(SADValues[790*12 +: 12], 12, 22, SADValues[727*12 +: 12], 11, 23, comp309minVal, comp309minI, comp309minJ);
    wire [11:0] comp310minVal;
    wire [5:0] comp310minI, comp310minJ;
    Comparator comp310(SADValues[664*12 +: 12], 10, 24, SADValues[601*12 +: 12], 9, 25, comp310minVal, comp310minI, comp310minJ);
    wire [11:0] comp311minVal;
    wire [5:0] comp311minI, comp311minJ;
    Comparator comp311(SADValues[538*12 +: 12], 8, 26, SADValues[475*12 +: 12], 7, 27, comp311minVal, comp311minI, comp311minJ);
    wire [11:0] comp312minVal;
    wire [5:0] comp312minI, comp312minJ;
    Comparator comp312(SADValues[412*12 +: 12], 6, 28, SADValues[349*12 +: 12], 5, 29, comp312minVal, comp312minI, comp312minJ);
    wire [11:0] comp313minVal;
    wire [5:0] comp313minI, comp313minJ;
    Comparator comp313(SADValues[286*12 +: 12], 4, 30, SADValues[223*12 +: 12], 3, 31, comp313minVal, comp313minI, comp313minJ);
    wire [11:0] comp314minVal;
    wire [5:0] comp314minI, comp314minJ;
    Comparator comp314(SADValues[160*12 +: 12], 2, 32, SADValues[97*12 +: 12], 1, 33, comp314minVal, comp314minI, comp314minJ);
    wire [11:0] comp315minVal;
    wire [5:0] comp315minI, comp315minJ;
    Comparator comp315(SADValues[34*12 +: 12], 0, 34, SADValues[35*12 +: 12], 0, 35, comp315minVal, comp315minI, comp315minJ);
    wire [11:0] comp316minVal;
    wire [5:0] comp316minI, comp316minJ;
    Comparator comp316(SADValues[98*12 +: 12], 1, 34, SADValues[161*12 +: 12], 2, 33, comp316minVal, comp316minI, comp316minJ);
    wire [11:0] comp317minVal;
    wire [5:0] comp317minI, comp317minJ;
    Comparator comp317(SADValues[224*12 +: 12], 3, 32, SADValues[287*12 +: 12], 4, 31, comp317minVal, comp317minI, comp317minJ);
    wire [11:0] comp318minVal;
    wire [5:0] comp318minI, comp318minJ;
    Comparator comp318(SADValues[350*12 +: 12], 5, 30, SADValues[413*12 +: 12], 6, 29, comp318minVal, comp318minI, comp318minJ);
    wire [11:0] comp319minVal;
    wire [5:0] comp319minI, comp319minJ;
    Comparator comp319(SADValues[476*12 +: 12], 7, 28, SADValues[539*12 +: 12], 8, 27, comp319minVal, comp319minI, comp319minJ);
    wire [11:0] comp320minVal;
    wire [5:0] comp320minI, comp320minJ;
    Comparator comp320(SADValues[602*12 +: 12], 9, 26, SADValues[665*12 +: 12], 10, 25, comp320minVal, comp320minI, comp320minJ);
    wire [11:0] comp321minVal;
    wire [5:0] comp321minI, comp321minJ;
    Comparator comp321(SADValues[728*12 +: 12], 11, 24, SADValues[791*12 +: 12], 12, 23, comp321minVal, comp321minI, comp321minJ);
    wire [11:0] comp322minVal;
    wire [5:0] comp322minI, comp322minJ;
    Comparator comp322(SADValues[854*12 +: 12], 13, 22, SADValues[917*12 +: 12], 14, 21, comp322minVal, comp322minI, comp322minJ);
    wire [11:0] comp323minVal;
    wire [5:0] comp323minI, comp323minJ;
    Comparator comp323(SADValues[980*12 +: 12], 15, 20, SADValues[1043*12 +: 12], 16, 19, comp323minVal, comp323minI, comp323minJ);
    wire [11:0] comp324minVal;
    wire [5:0] comp324minI, comp324minJ;
    Comparator comp324(SADValues[1106*12 +: 12], 17, 18, SADValues[1169*12 +: 12], 18, 17, comp324minVal, comp324minI, comp324minJ);
    wire [11:0] comp325minVal;
    wire [5:0] comp325minI, comp325minJ;
    Comparator comp325(SADValues[1232*12 +: 12], 19, 16, SADValues[1295*12 +: 12], 20, 15, comp325minVal, comp325minI, comp325minJ);
    wire [11:0] comp326minVal;
    wire [5:0] comp326minI, comp326minJ;
    Comparator comp326(SADValues[1358*12 +: 12], 21, 14, SADValues[1421*12 +: 12], 22, 13, comp326minVal, comp326minI, comp326minJ);
    wire [11:0] comp327minVal;
    wire [5:0] comp327minI, comp327minJ;
    Comparator comp327(SADValues[1484*12 +: 12], 23, 12, SADValues[1547*12 +: 12], 24, 11, comp327minVal, comp327minI, comp327minJ);
    wire [11:0] comp328minVal;
    wire [5:0] comp328minI, comp328minJ;
    Comparator comp328(SADValues[1610*12 +: 12], 25, 10, SADValues[1673*12 +: 12], 26, 9, comp328minVal, comp328minI, comp328minJ);
    wire [11:0] comp329minVal;
    wire [5:0] comp329minI, comp329minJ;
    Comparator comp329(SADValues[1736*12 +: 12], 27, 8, SADValues[1799*12 +: 12], 28, 7, comp329minVal, comp329minI, comp329minJ);
    wire [11:0] comp330minVal;
    wire [5:0] comp330minI, comp330minJ;
    Comparator comp330(SADValues[1862*12 +: 12], 29, 6, SADValues[1925*12 +: 12], 30, 5, comp330minVal, comp330minI, comp330minJ);
    wire [11:0] comp331minVal;
    wire [5:0] comp331minI, comp331minJ;
    Comparator comp331(SADValues[1988*12 +: 12], 31, 4, SADValues[2051*12 +: 12], 32, 3, comp331minVal, comp331minI, comp331minJ);
    wire [11:0] comp332minVal;
    wire [5:0] comp332minI, comp332minJ;
    Comparator comp332(SADValues[2114*12 +: 12], 33, 2, SADValues[2177*12 +: 12], 34, 1, comp332minVal, comp332minI, comp332minJ);
    wire [11:0] comp333minVal;
    wire [5:0] comp333minI, comp333minJ;
    Comparator comp333(SADValues[2240*12 +: 12], 35, 0, SADValues[2304*12 +: 12], 36, 0, comp333minVal, comp333minI, comp333minJ);
    wire [11:0] comp334minVal;
    wire [5:0] comp334minI, comp334minJ;
    Comparator comp334(SADValues[2241*12 +: 12], 35, 1, SADValues[2178*12 +: 12], 34, 2, comp334minVal, comp334minI, comp334minJ);
    wire [11:0] comp335minVal;
    wire [5:0] comp335minI, comp335minJ;
    Comparator comp335(SADValues[2115*12 +: 12], 33, 3, SADValues[2052*12 +: 12], 32, 4, comp335minVal, comp335minI, comp335minJ);
    wire [11:0] comp336minVal;
    wire [5:0] comp336minI, comp336minJ;
    Comparator comp336(SADValues[1989*12 +: 12], 31, 5, SADValues[1926*12 +: 12], 30, 6, comp336minVal, comp336minI, comp336minJ);
    wire [11:0] comp337minVal;
    wire [5:0] comp337minI, comp337minJ;
    Comparator comp337(SADValues[1863*12 +: 12], 29, 7, SADValues[1800*12 +: 12], 28, 8, comp337minVal, comp337minI, comp337minJ);
    wire [11:0] comp338minVal;
    wire [5:0] comp338minI, comp338minJ;
    Comparator comp338(SADValues[1737*12 +: 12], 27, 9, SADValues[1674*12 +: 12], 26, 10, comp338minVal, comp338minI, comp338minJ);
    wire [11:0] comp339minVal;
    wire [5:0] comp339minI, comp339minJ;
    Comparator comp339(SADValues[1611*12 +: 12], 25, 11, SADValues[1548*12 +: 12], 24, 12, comp339minVal, comp339minI, comp339minJ);
    wire [11:0] comp340minVal;
    wire [5:0] comp340minI, comp340minJ;
    Comparator comp340(SADValues[1485*12 +: 12], 23, 13, SADValues[1422*12 +: 12], 22, 14, comp340minVal, comp340minI, comp340minJ);
    wire [11:0] comp341minVal;
    wire [5:0] comp341minI, comp341minJ;
    Comparator comp341(SADValues[1359*12 +: 12], 21, 15, SADValues[1296*12 +: 12], 20, 16, comp341minVal, comp341minI, comp341minJ);
    wire [11:0] comp342minVal;
    wire [5:0] comp342minI, comp342minJ;
    Comparator comp342(SADValues[1233*12 +: 12], 19, 17, SADValues[1170*12 +: 12], 18, 18, comp342minVal, comp342minI, comp342minJ);
    wire [11:0] comp343minVal;
    wire [5:0] comp343minI, comp343minJ;
    Comparator comp343(SADValues[1107*12 +: 12], 17, 19, SADValues[1044*12 +: 12], 16, 20, comp343minVal, comp343minI, comp343minJ);
    wire [11:0] comp344minVal;
    wire [5:0] comp344minI, comp344minJ;
    Comparator comp344(SADValues[981*12 +: 12], 15, 21, SADValues[918*12 +: 12], 14, 22, comp344minVal, comp344minI, comp344minJ);
    wire [11:0] comp345minVal;
    wire [5:0] comp345minI, comp345minJ;
    Comparator comp345(SADValues[855*12 +: 12], 13, 23, SADValues[792*12 +: 12], 12, 24, comp345minVal, comp345minI, comp345minJ);
    wire [11:0] comp346minVal;
    wire [5:0] comp346minI, comp346minJ;
    Comparator comp346(SADValues[729*12 +: 12], 11, 25, SADValues[666*12 +: 12], 10, 26, comp346minVal, comp346minI, comp346minJ);
    wire [11:0] comp347minVal;
    wire [5:0] comp347minI, comp347minJ;
    Comparator comp347(SADValues[603*12 +: 12], 9, 27, SADValues[540*12 +: 12], 8, 28, comp347minVal, comp347minI, comp347minJ);
    wire [11:0] comp348minVal;
    wire [5:0] comp348minI, comp348minJ;
    Comparator comp348(SADValues[477*12 +: 12], 7, 29, SADValues[414*12 +: 12], 6, 30, comp348minVal, comp348minI, comp348minJ);
    wire [11:0] comp349minVal;
    wire [5:0] comp349minI, comp349minJ;
    Comparator comp349(SADValues[351*12 +: 12], 5, 31, SADValues[288*12 +: 12], 4, 32, comp349minVal, comp349minI, comp349minJ);
    wire [11:0] comp350minVal;
    wire [5:0] comp350minI, comp350minJ;
    Comparator comp350(SADValues[225*12 +: 12], 3, 33, SADValues[162*12 +: 12], 2, 34, comp350minVal, comp350minI, comp350minJ);
    wire [11:0] comp351minVal;
    wire [5:0] comp351minI, comp351minJ;
    Comparator comp351(SADValues[99*12 +: 12], 1, 35, SADValues[36*12 +: 12], 0, 36, comp351minVal, comp351minI, comp351minJ);
    wire [11:0] comp352minVal;
    wire [5:0] comp352minI, comp352minJ;
    Comparator comp352(SADValues[37*12 +: 12], 0, 37, SADValues[100*12 +: 12], 1, 36, comp352minVal, comp352minI, comp352minJ);
    wire [11:0] comp353minVal;
    wire [5:0] comp353minI, comp353minJ;
    Comparator comp353(SADValues[163*12 +: 12], 2, 35, SADValues[226*12 +: 12], 3, 34, comp353minVal, comp353minI, comp353minJ);
    wire [11:0] comp354minVal;
    wire [5:0] comp354minI, comp354minJ;
    Comparator comp354(SADValues[289*12 +: 12], 4, 33, SADValues[352*12 +: 12], 5, 32, comp354minVal, comp354minI, comp354minJ);
    wire [11:0] comp355minVal;
    wire [5:0] comp355minI, comp355minJ;
    Comparator comp355(SADValues[415*12 +: 12], 6, 31, SADValues[478*12 +: 12], 7, 30, comp355minVal, comp355minI, comp355minJ);
    wire [11:0] comp356minVal;
    wire [5:0] comp356minI, comp356minJ;
    Comparator comp356(SADValues[541*12 +: 12], 8, 29, SADValues[604*12 +: 12], 9, 28, comp356minVal, comp356minI, comp356minJ);
    wire [11:0] comp357minVal;
    wire [5:0] comp357minI, comp357minJ;
    Comparator comp357(SADValues[667*12 +: 12], 10, 27, SADValues[730*12 +: 12], 11, 26, comp357minVal, comp357minI, comp357minJ);
    wire [11:0] comp358minVal;
    wire [5:0] comp358minI, comp358minJ;
    Comparator comp358(SADValues[793*12 +: 12], 12, 25, SADValues[856*12 +: 12], 13, 24, comp358minVal, comp358minI, comp358minJ);
    wire [11:0] comp359minVal;
    wire [5:0] comp359minI, comp359minJ;
    Comparator comp359(SADValues[919*12 +: 12], 14, 23, SADValues[982*12 +: 12], 15, 22, comp359minVal, comp359minI, comp359minJ);
    wire [11:0] comp360minVal;
    wire [5:0] comp360minI, comp360minJ;
    Comparator comp360(SADValues[1045*12 +: 12], 16, 21, SADValues[1108*12 +: 12], 17, 20, comp360minVal, comp360minI, comp360minJ);
    wire [11:0] comp361minVal;
    wire [5:0] comp361minI, comp361minJ;
    Comparator comp361(SADValues[1171*12 +: 12], 18, 19, SADValues[1234*12 +: 12], 19, 18, comp361minVal, comp361minI, comp361minJ);
    wire [11:0] comp362minVal;
    wire [5:0] comp362minI, comp362minJ;
    Comparator comp362(SADValues[1297*12 +: 12], 20, 17, SADValues[1360*12 +: 12], 21, 16, comp362minVal, comp362minI, comp362minJ);
    wire [11:0] comp363minVal;
    wire [5:0] comp363minI, comp363minJ;
    Comparator comp363(SADValues[1423*12 +: 12], 22, 15, SADValues[1486*12 +: 12], 23, 14, comp363minVal, comp363minI, comp363minJ);
    wire [11:0] comp364minVal;
    wire [5:0] comp364minI, comp364minJ;
    Comparator comp364(SADValues[1549*12 +: 12], 24, 13, SADValues[1612*12 +: 12], 25, 12, comp364minVal, comp364minI, comp364minJ);
    wire [11:0] comp365minVal;
    wire [5:0] comp365minI, comp365minJ;
    Comparator comp365(SADValues[1675*12 +: 12], 26, 11, SADValues[1738*12 +: 12], 27, 10, comp365minVal, comp365minI, comp365minJ);
    wire [11:0] comp366minVal;
    wire [5:0] comp366minI, comp366minJ;
    Comparator comp366(SADValues[1801*12 +: 12], 28, 9, SADValues[1864*12 +: 12], 29, 8, comp366minVal, comp366minI, comp366minJ);
    wire [11:0] comp367minVal;
    wire [5:0] comp367minI, comp367minJ;
    Comparator comp367(SADValues[1927*12 +: 12], 30, 7, SADValues[1990*12 +: 12], 31, 6, comp367minVal, comp367minI, comp367minJ);
    wire [11:0] comp368minVal;
    wire [5:0] comp368minI, comp368minJ;
    Comparator comp368(SADValues[2053*12 +: 12], 32, 5, SADValues[2116*12 +: 12], 33, 4, comp368minVal, comp368minI, comp368minJ);
    wire [11:0] comp369minVal;
    wire [5:0] comp369minI, comp369minJ;
    Comparator comp369(SADValues[2179*12 +: 12], 34, 3, SADValues[2242*12 +: 12], 35, 2, comp369minVal, comp369minI, comp369minJ);
    wire [11:0] comp370minVal;
    wire [5:0] comp370minI, comp370minJ;
    Comparator comp370(SADValues[2305*12 +: 12], 36, 1, SADValues[2368*12 +: 12], 37, 0, comp370minVal, comp370minI, comp370minJ);
    wire [11:0] comp371minVal;
    wire [5:0] comp371minI, comp371minJ;
    Comparator comp371(SADValues[2432*12 +: 12], 38, 0, SADValues[2369*12 +: 12], 37, 1, comp371minVal, comp371minI, comp371minJ);
    wire [11:0] comp372minVal;
    wire [5:0] comp372minI, comp372minJ;
    Comparator comp372(SADValues[2306*12 +: 12], 36, 2, SADValues[2243*12 +: 12], 35, 3, comp372minVal, comp372minI, comp372minJ);
    wire [11:0] comp373minVal;
    wire [5:0] comp373minI, comp373minJ;
    Comparator comp373(SADValues[2180*12 +: 12], 34, 4, SADValues[2117*12 +: 12], 33, 5, comp373minVal, comp373minI, comp373minJ);
    wire [11:0] comp374minVal;
    wire [5:0] comp374minI, comp374minJ;
    Comparator comp374(SADValues[2054*12 +: 12], 32, 6, SADValues[1991*12 +: 12], 31, 7, comp374minVal, comp374minI, comp374minJ);
    wire [11:0] comp375minVal;
    wire [5:0] comp375minI, comp375minJ;
    Comparator comp375(SADValues[1928*12 +: 12], 30, 8, SADValues[1865*12 +: 12], 29, 9, comp375minVal, comp375minI, comp375minJ);
    wire [11:0] comp376minVal;
    wire [5:0] comp376minI, comp376minJ;
    Comparator comp376(SADValues[1802*12 +: 12], 28, 10, SADValues[1739*12 +: 12], 27, 11, comp376minVal, comp376minI, comp376minJ);
    wire [11:0] comp377minVal;
    wire [5:0] comp377minI, comp377minJ;
    Comparator comp377(SADValues[1676*12 +: 12], 26, 12, SADValues[1613*12 +: 12], 25, 13, comp377minVal, comp377minI, comp377minJ);
    wire [11:0] comp378minVal;
    wire [5:0] comp378minI, comp378minJ;
    Comparator comp378(SADValues[1550*12 +: 12], 24, 14, SADValues[1487*12 +: 12], 23, 15, comp378minVal, comp378minI, comp378minJ);
    wire [11:0] comp379minVal;
    wire [5:0] comp379minI, comp379minJ;
    Comparator comp379(SADValues[1424*12 +: 12], 22, 16, SADValues[1361*12 +: 12], 21, 17, comp379minVal, comp379minI, comp379minJ);
    wire [11:0] comp380minVal;
    wire [5:0] comp380minI, comp380minJ;
    Comparator comp380(SADValues[1298*12 +: 12], 20, 18, SADValues[1235*12 +: 12], 19, 19, comp380minVal, comp380minI, comp380minJ);
    wire [11:0] comp381minVal;
    wire [5:0] comp381minI, comp381minJ;
    Comparator comp381(SADValues[1172*12 +: 12], 18, 20, SADValues[1109*12 +: 12], 17, 21, comp381minVal, comp381minI, comp381minJ);
    wire [11:0] comp382minVal;
    wire [5:0] comp382minI, comp382minJ;
    Comparator comp382(SADValues[1046*12 +: 12], 16, 22, SADValues[983*12 +: 12], 15, 23, comp382minVal, comp382minI, comp382minJ);
    wire [11:0] comp383minVal;
    wire [5:0] comp383minI, comp383minJ;
    Comparator comp383(SADValues[920*12 +: 12], 14, 24, SADValues[857*12 +: 12], 13, 25, comp383minVal, comp383minI, comp383minJ);
    wire [11:0] comp384minVal;
    wire [5:0] comp384minI, comp384minJ;
    Comparator comp384(SADValues[794*12 +: 12], 12, 26, SADValues[731*12 +: 12], 11, 27, comp384minVal, comp384minI, comp384minJ);
    wire [11:0] comp385minVal;
    wire [5:0] comp385minI, comp385minJ;
    Comparator comp385(SADValues[668*12 +: 12], 10, 28, SADValues[605*12 +: 12], 9, 29, comp385minVal, comp385minI, comp385minJ);
    wire [11:0] comp386minVal;
    wire [5:0] comp386minI, comp386minJ;
    Comparator comp386(SADValues[542*12 +: 12], 8, 30, SADValues[479*12 +: 12], 7, 31, comp386minVal, comp386minI, comp386minJ);
    wire [11:0] comp387minVal;
    wire [5:0] comp387minI, comp387minJ;
    Comparator comp387(SADValues[416*12 +: 12], 6, 32, SADValues[353*12 +: 12], 5, 33, comp387minVal, comp387minI, comp387minJ);
    wire [11:0] comp388minVal;
    wire [5:0] comp388minI, comp388minJ;
    Comparator comp388(SADValues[290*12 +: 12], 4, 34, SADValues[227*12 +: 12], 3, 35, comp388minVal, comp388minI, comp388minJ);
    wire [11:0] comp389minVal;
    wire [5:0] comp389minI, comp389minJ;
    Comparator comp389(SADValues[164*12 +: 12], 2, 36, SADValues[101*12 +: 12], 1, 37, comp389minVal, comp389minI, comp389minJ);
    wire [11:0] comp390minVal;
    wire [5:0] comp390minI, comp390minJ;
    Comparator comp390(SADValues[38*12 +: 12], 0, 38, SADValues[39*12 +: 12], 0, 39, comp390minVal, comp390minI, comp390minJ);
    wire [11:0] comp391minVal;
    wire [5:0] comp391minI, comp391minJ;
    Comparator comp391(SADValues[102*12 +: 12], 1, 38, SADValues[165*12 +: 12], 2, 37, comp391minVal, comp391minI, comp391minJ);
    wire [11:0] comp392minVal;
    wire [5:0] comp392minI, comp392minJ;
    Comparator comp392(SADValues[228*12 +: 12], 3, 36, SADValues[291*12 +: 12], 4, 35, comp392minVal, comp392minI, comp392minJ);
    wire [11:0] comp393minVal;
    wire [5:0] comp393minI, comp393minJ;
    Comparator comp393(SADValues[354*12 +: 12], 5, 34, SADValues[417*12 +: 12], 6, 33, comp393minVal, comp393minI, comp393minJ);
    wire [11:0] comp394minVal;
    wire [5:0] comp394minI, comp394minJ;
    Comparator comp394(SADValues[480*12 +: 12], 7, 32, SADValues[543*12 +: 12], 8, 31, comp394minVal, comp394minI, comp394minJ);
    wire [11:0] comp395minVal;
    wire [5:0] comp395minI, comp395minJ;
    Comparator comp395(SADValues[606*12 +: 12], 9, 30, SADValues[669*12 +: 12], 10, 29, comp395minVal, comp395minI, comp395minJ);
    wire [11:0] comp396minVal;
    wire [5:0] comp396minI, comp396minJ;
    Comparator comp396(SADValues[732*12 +: 12], 11, 28, SADValues[795*12 +: 12], 12, 27, comp396minVal, comp396minI, comp396minJ);
    wire [11:0] comp397minVal;
    wire [5:0] comp397minI, comp397minJ;
    Comparator comp397(SADValues[858*12 +: 12], 13, 26, SADValues[921*12 +: 12], 14, 25, comp397minVal, comp397minI, comp397minJ);
    wire [11:0] comp398minVal;
    wire [5:0] comp398minI, comp398minJ;
    Comparator comp398(SADValues[984*12 +: 12], 15, 24, SADValues[1047*12 +: 12], 16, 23, comp398minVal, comp398minI, comp398minJ);
    wire [11:0] comp399minVal;
    wire [5:0] comp399minI, comp399minJ;
    Comparator comp399(SADValues[1110*12 +: 12], 17, 22, SADValues[1173*12 +: 12], 18, 21, comp399minVal, comp399minI, comp399minJ);
    wire [11:0] comp400minVal;
    wire [5:0] comp400minI, comp400minJ;
    Comparator comp400(SADValues[1236*12 +: 12], 19, 20, SADValues[1299*12 +: 12], 20, 19, comp400minVal, comp400minI, comp400minJ);
    wire [11:0] comp401minVal;
    wire [5:0] comp401minI, comp401minJ;
    Comparator comp401(SADValues[1362*12 +: 12], 21, 18, SADValues[1425*12 +: 12], 22, 17, comp401minVal, comp401minI, comp401minJ);
    wire [11:0] comp402minVal;
    wire [5:0] comp402minI, comp402minJ;
    Comparator comp402(SADValues[1488*12 +: 12], 23, 16, SADValues[1551*12 +: 12], 24, 15, comp402minVal, comp402minI, comp402minJ);
    wire [11:0] comp403minVal;
    wire [5:0] comp403minI, comp403minJ;
    Comparator comp403(SADValues[1614*12 +: 12], 25, 14, SADValues[1677*12 +: 12], 26, 13, comp403minVal, comp403minI, comp403minJ);
    wire [11:0] comp404minVal;
    wire [5:0] comp404minI, comp404minJ;
    Comparator comp404(SADValues[1740*12 +: 12], 27, 12, SADValues[1803*12 +: 12], 28, 11, comp404minVal, comp404minI, comp404minJ);
    wire [11:0] comp405minVal;
    wire [5:0] comp405minI, comp405minJ;
    Comparator comp405(SADValues[1866*12 +: 12], 29, 10, SADValues[1929*12 +: 12], 30, 9, comp405minVal, comp405minI, comp405minJ);
    wire [11:0] comp406minVal;
    wire [5:0] comp406minI, comp406minJ;
    Comparator comp406(SADValues[1992*12 +: 12], 31, 8, SADValues[2055*12 +: 12], 32, 7, comp406minVal, comp406minI, comp406minJ);
    wire [11:0] comp407minVal;
    wire [5:0] comp407minI, comp407minJ;
    Comparator comp407(SADValues[2118*12 +: 12], 33, 6, SADValues[2181*12 +: 12], 34, 5, comp407minVal, comp407minI, comp407minJ);
    wire [11:0] comp408minVal;
    wire [5:0] comp408minI, comp408minJ;
    Comparator comp408(SADValues[2244*12 +: 12], 35, 4, SADValues[2307*12 +: 12], 36, 3, comp408minVal, comp408minI, comp408minJ);
    wire [11:0] comp409minVal;
    wire [5:0] comp409minI, comp409minJ;
    Comparator comp409(SADValues[2370*12 +: 12], 37, 2, SADValues[2433*12 +: 12], 38, 1, comp409minVal, comp409minI, comp409minJ);
    wire [11:0] comp410minVal;
    wire [5:0] comp410minI, comp410minJ;
    Comparator comp410(SADValues[2496*12 +: 12], 39, 0, SADValues[2560*12 +: 12], 40, 0, comp410minVal, comp410minI, comp410minJ);
    wire [11:0] comp411minVal;
    wire [5:0] comp411minI, comp411minJ;
    Comparator comp411(SADValues[2497*12 +: 12], 39, 1, SADValues[2434*12 +: 12], 38, 2, comp411minVal, comp411minI, comp411minJ);
    wire [11:0] comp412minVal;
    wire [5:0] comp412minI, comp412minJ;
    Comparator comp412(SADValues[2371*12 +: 12], 37, 3, SADValues[2308*12 +: 12], 36, 4, comp412minVal, comp412minI, comp412minJ);
    wire [11:0] comp413minVal;
    wire [5:0] comp413minI, comp413minJ;
    Comparator comp413(SADValues[2245*12 +: 12], 35, 5, SADValues[2182*12 +: 12], 34, 6, comp413minVal, comp413minI, comp413minJ);
    wire [11:0] comp414minVal;
    wire [5:0] comp414minI, comp414minJ;
    Comparator comp414(SADValues[2119*12 +: 12], 33, 7, SADValues[2056*12 +: 12], 32, 8, comp414minVal, comp414minI, comp414minJ);
    wire [11:0] comp415minVal;
    wire [5:0] comp415minI, comp415minJ;
    Comparator comp415(SADValues[1993*12 +: 12], 31, 9, SADValues[1930*12 +: 12], 30, 10, comp415minVal, comp415minI, comp415minJ);
    wire [11:0] comp416minVal;
    wire [5:0] comp416minI, comp416minJ;
    Comparator comp416(SADValues[1867*12 +: 12], 29, 11, SADValues[1804*12 +: 12], 28, 12, comp416minVal, comp416minI, comp416minJ);
    wire [11:0] comp417minVal;
    wire [5:0] comp417minI, comp417minJ;
    Comparator comp417(SADValues[1741*12 +: 12], 27, 13, SADValues[1678*12 +: 12], 26, 14, comp417minVal, comp417minI, comp417minJ);
    wire [11:0] comp418minVal;
    wire [5:0] comp418minI, comp418minJ;
    Comparator comp418(SADValues[1615*12 +: 12], 25, 15, SADValues[1552*12 +: 12], 24, 16, comp418minVal, comp418minI, comp418minJ);
    wire [11:0] comp419minVal;
    wire [5:0] comp419minI, comp419minJ;
    Comparator comp419(SADValues[1489*12 +: 12], 23, 17, SADValues[1426*12 +: 12], 22, 18, comp419minVal, comp419minI, comp419minJ);
    wire [11:0] comp420minVal;
    wire [5:0] comp420minI, comp420minJ;
    Comparator comp420(SADValues[1363*12 +: 12], 21, 19, SADValues[1300*12 +: 12], 20, 20, comp420minVal, comp420minI, comp420minJ);
    wire [11:0] comp421minVal;
    wire [5:0] comp421minI, comp421minJ;
    Comparator comp421(SADValues[1237*12 +: 12], 19, 21, SADValues[1174*12 +: 12], 18, 22, comp421minVal, comp421minI, comp421minJ);
    wire [11:0] comp422minVal;
    wire [5:0] comp422minI, comp422minJ;
    Comparator comp422(SADValues[1111*12 +: 12], 17, 23, SADValues[1048*12 +: 12], 16, 24, comp422minVal, comp422minI, comp422minJ);
    wire [11:0] comp423minVal;
    wire [5:0] comp423minI, comp423minJ;
    Comparator comp423(SADValues[985*12 +: 12], 15, 25, SADValues[922*12 +: 12], 14, 26, comp423minVal, comp423minI, comp423minJ);
    wire [11:0] comp424minVal;
    wire [5:0] comp424minI, comp424minJ;
    Comparator comp424(SADValues[859*12 +: 12], 13, 27, SADValues[796*12 +: 12], 12, 28, comp424minVal, comp424minI, comp424minJ);
    wire [11:0] comp425minVal;
    wire [5:0] comp425minI, comp425minJ;
    Comparator comp425(SADValues[733*12 +: 12], 11, 29, SADValues[670*12 +: 12], 10, 30, comp425minVal, comp425minI, comp425minJ);
    wire [11:0] comp426minVal;
    wire [5:0] comp426minI, comp426minJ;
    Comparator comp426(SADValues[607*12 +: 12], 9, 31, SADValues[544*12 +: 12], 8, 32, comp426minVal, comp426minI, comp426minJ);
    wire [11:0] comp427minVal;
    wire [5:0] comp427minI, comp427minJ;
    Comparator comp427(SADValues[481*12 +: 12], 7, 33, SADValues[418*12 +: 12], 6, 34, comp427minVal, comp427minI, comp427minJ);
    wire [11:0] comp428minVal;
    wire [5:0] comp428minI, comp428minJ;
    Comparator comp428(SADValues[355*12 +: 12], 5, 35, SADValues[292*12 +: 12], 4, 36, comp428minVal, comp428minI, comp428minJ);
    wire [11:0] comp429minVal;
    wire [5:0] comp429minI, comp429minJ;
    Comparator comp429(SADValues[229*12 +: 12], 3, 37, SADValues[166*12 +: 12], 2, 38, comp429minVal, comp429minI, comp429minJ);
    wire [11:0] comp430minVal;
    wire [5:0] comp430minI, comp430minJ;
    Comparator comp430(SADValues[103*12 +: 12], 1, 39, SADValues[40*12 +: 12], 0, 40, comp430minVal, comp430minI, comp430minJ);
    wire [11:0] comp431minVal;
    wire [5:0] comp431minI, comp431minJ;
    Comparator comp431(SADValues[41*12 +: 12], 0, 41, SADValues[104*12 +: 12], 1, 40, comp431minVal, comp431minI, comp431minJ);
    wire [11:0] comp432minVal;
    wire [5:0] comp432minI, comp432minJ;
    Comparator comp432(SADValues[167*12 +: 12], 2, 39, SADValues[230*12 +: 12], 3, 38, comp432minVal, comp432minI, comp432minJ);
    wire [11:0] comp433minVal;
    wire [5:0] comp433minI, comp433minJ;
    Comparator comp433(SADValues[293*12 +: 12], 4, 37, SADValues[356*12 +: 12], 5, 36, comp433minVal, comp433minI, comp433minJ);
    wire [11:0] comp434minVal;
    wire [5:0] comp434minI, comp434minJ;
    Comparator comp434(SADValues[419*12 +: 12], 6, 35, SADValues[482*12 +: 12], 7, 34, comp434minVal, comp434minI, comp434minJ);
    wire [11:0] comp435minVal;
    wire [5:0] comp435minI, comp435minJ;
    Comparator comp435(SADValues[545*12 +: 12], 8, 33, SADValues[608*12 +: 12], 9, 32, comp435minVal, comp435minI, comp435minJ);
    wire [11:0] comp436minVal;
    wire [5:0] comp436minI, comp436minJ;
    Comparator comp436(SADValues[671*12 +: 12], 10, 31, SADValues[734*12 +: 12], 11, 30, comp436minVal, comp436minI, comp436minJ);
    wire [11:0] comp437minVal;
    wire [5:0] comp437minI, comp437minJ;
    Comparator comp437(SADValues[797*12 +: 12], 12, 29, SADValues[860*12 +: 12], 13, 28, comp437minVal, comp437minI, comp437minJ);
    wire [11:0] comp438minVal;
    wire [5:0] comp438minI, comp438minJ;
    Comparator comp438(SADValues[923*12 +: 12], 14, 27, SADValues[986*12 +: 12], 15, 26, comp438minVal, comp438minI, comp438minJ);
    wire [11:0] comp439minVal;
    wire [5:0] comp439minI, comp439minJ;
    Comparator comp439(SADValues[1049*12 +: 12], 16, 25, SADValues[1112*12 +: 12], 17, 24, comp439minVal, comp439minI, comp439minJ);
    wire [11:0] comp440minVal;
    wire [5:0] comp440minI, comp440minJ;
    Comparator comp440(SADValues[1175*12 +: 12], 18, 23, SADValues[1238*12 +: 12], 19, 22, comp440minVal, comp440minI, comp440minJ);
    wire [11:0] comp441minVal;
    wire [5:0] comp441minI, comp441minJ;
    Comparator comp441(SADValues[1301*12 +: 12], 20, 21, SADValues[1364*12 +: 12], 21, 20, comp441minVal, comp441minI, comp441minJ);
    wire [11:0] comp442minVal;
    wire [5:0] comp442minI, comp442minJ;
    Comparator comp442(SADValues[1427*12 +: 12], 22, 19, SADValues[1490*12 +: 12], 23, 18, comp442minVal, comp442minI, comp442minJ);
    wire [11:0] comp443minVal;
    wire [5:0] comp443minI, comp443minJ;
    Comparator comp443(SADValues[1553*12 +: 12], 24, 17, SADValues[1616*12 +: 12], 25, 16, comp443minVal, comp443minI, comp443minJ);
    wire [11:0] comp444minVal;
    wire [5:0] comp444minI, comp444minJ;
    Comparator comp444(SADValues[1679*12 +: 12], 26, 15, SADValues[1742*12 +: 12], 27, 14, comp444minVal, comp444minI, comp444minJ);
    wire [11:0] comp445minVal;
    wire [5:0] comp445minI, comp445minJ;
    Comparator comp445(SADValues[1805*12 +: 12], 28, 13, SADValues[1868*12 +: 12], 29, 12, comp445minVal, comp445minI, comp445minJ);
    wire [11:0] comp446minVal;
    wire [5:0] comp446minI, comp446minJ;
    Comparator comp446(SADValues[1931*12 +: 12], 30, 11, SADValues[1994*12 +: 12], 31, 10, comp446minVal, comp446minI, comp446minJ);
    wire [11:0] comp447minVal;
    wire [5:0] comp447minI, comp447minJ;
    Comparator comp447(SADValues[2057*12 +: 12], 32, 9, SADValues[2120*12 +: 12], 33, 8, comp447minVal, comp447minI, comp447minJ);
    wire [11:0] comp448minVal;
    wire [5:0] comp448minI, comp448minJ;
    Comparator comp448(SADValues[2183*12 +: 12], 34, 7, SADValues[2246*12 +: 12], 35, 6, comp448minVal, comp448minI, comp448minJ);
    wire [11:0] comp449minVal;
    wire [5:0] comp449minI, comp449minJ;
    Comparator comp449(SADValues[2309*12 +: 12], 36, 5, SADValues[2372*12 +: 12], 37, 4, comp449minVal, comp449minI, comp449minJ);
    wire [11:0] comp450minVal;
    wire [5:0] comp450minI, comp450minJ;
    Comparator comp450(SADValues[2435*12 +: 12], 38, 3, SADValues[2498*12 +: 12], 39, 2, comp450minVal, comp450minI, comp450minJ);
    wire [11:0] comp451minVal;
    wire [5:0] comp451minI, comp451minJ;
    Comparator comp451(SADValues[2561*12 +: 12], 40, 1, SADValues[2624*12 +: 12], 41, 0, comp451minVal, comp451minI, comp451minJ);
    wire [11:0] comp452minVal;
    wire [5:0] comp452minI, comp452minJ;
    Comparator comp452(SADValues[2688*12 +: 12], 42, 0, SADValues[2625*12 +: 12], 41, 1, comp452minVal, comp452minI, comp452minJ);
    wire [11:0] comp453minVal;
    wire [5:0] comp453minI, comp453minJ;
    Comparator comp453(SADValues[2562*12 +: 12], 40, 2, SADValues[2499*12 +: 12], 39, 3, comp453minVal, comp453minI, comp453minJ);
    wire [11:0] comp454minVal;
    wire [5:0] comp454minI, comp454minJ;
    Comparator comp454(SADValues[2436*12 +: 12], 38, 4, SADValues[2373*12 +: 12], 37, 5, comp454minVal, comp454minI, comp454minJ);
    wire [11:0] comp455minVal;
    wire [5:0] comp455minI, comp455minJ;
    Comparator comp455(SADValues[2310*12 +: 12], 36, 6, SADValues[2247*12 +: 12], 35, 7, comp455minVal, comp455minI, comp455minJ);
    wire [11:0] comp456minVal;
    wire [5:0] comp456minI, comp456minJ;
    Comparator comp456(SADValues[2184*12 +: 12], 34, 8, SADValues[2121*12 +: 12], 33, 9, comp456minVal, comp456minI, comp456minJ);
    wire [11:0] comp457minVal;
    wire [5:0] comp457minI, comp457minJ;
    Comparator comp457(SADValues[2058*12 +: 12], 32, 10, SADValues[1995*12 +: 12], 31, 11, comp457minVal, comp457minI, comp457minJ);
    wire [11:0] comp458minVal;
    wire [5:0] comp458minI, comp458minJ;
    Comparator comp458(SADValues[1932*12 +: 12], 30, 12, SADValues[1869*12 +: 12], 29, 13, comp458minVal, comp458minI, comp458minJ);
    wire [11:0] comp459minVal;
    wire [5:0] comp459minI, comp459minJ;
    Comparator comp459(SADValues[1806*12 +: 12], 28, 14, SADValues[1743*12 +: 12], 27, 15, comp459minVal, comp459minI, comp459minJ);
    wire [11:0] comp460minVal;
    wire [5:0] comp460minI, comp460minJ;
    Comparator comp460(SADValues[1680*12 +: 12], 26, 16, SADValues[1617*12 +: 12], 25, 17, comp460minVal, comp460minI, comp460minJ);
    wire [11:0] comp461minVal;
    wire [5:0] comp461minI, comp461minJ;
    Comparator comp461(SADValues[1554*12 +: 12], 24, 18, SADValues[1491*12 +: 12], 23, 19, comp461minVal, comp461minI, comp461minJ);
    wire [11:0] comp462minVal;
    wire [5:0] comp462minI, comp462minJ;
    Comparator comp462(SADValues[1428*12 +: 12], 22, 20, SADValues[1365*12 +: 12], 21, 21, comp462minVal, comp462minI, comp462minJ);
    wire [11:0] comp463minVal;
    wire [5:0] comp463minI, comp463minJ;
    Comparator comp463(SADValues[1302*12 +: 12], 20, 22, SADValues[1239*12 +: 12], 19, 23, comp463minVal, comp463minI, comp463minJ);
    wire [11:0] comp464minVal;
    wire [5:0] comp464minI, comp464minJ;
    Comparator comp464(SADValues[1176*12 +: 12], 18, 24, SADValues[1113*12 +: 12], 17, 25, comp464minVal, comp464minI, comp464minJ);
    wire [11:0] comp465minVal;
    wire [5:0] comp465minI, comp465minJ;
    Comparator comp465(SADValues[1050*12 +: 12], 16, 26, SADValues[987*12 +: 12], 15, 27, comp465minVal, comp465minI, comp465minJ);
    wire [11:0] comp466minVal;
    wire [5:0] comp466minI, comp466minJ;
    Comparator comp466(SADValues[924*12 +: 12], 14, 28, SADValues[861*12 +: 12], 13, 29, comp466minVal, comp466minI, comp466minJ);
    wire [11:0] comp467minVal;
    wire [5:0] comp467minI, comp467minJ;
    Comparator comp467(SADValues[798*12 +: 12], 12, 30, SADValues[735*12 +: 12], 11, 31, comp467minVal, comp467minI, comp467minJ);
    wire [11:0] comp468minVal;
    wire [5:0] comp468minI, comp468minJ;
    Comparator comp468(SADValues[672*12 +: 12], 10, 32, SADValues[609*12 +: 12], 9, 33, comp468minVal, comp468minI, comp468minJ);
    wire [11:0] comp469minVal;
    wire [5:0] comp469minI, comp469minJ;
    Comparator comp469(SADValues[546*12 +: 12], 8, 34, SADValues[483*12 +: 12], 7, 35, comp469minVal, comp469minI, comp469minJ);
    wire [11:0] comp470minVal;
    wire [5:0] comp470minI, comp470minJ;
    Comparator comp470(SADValues[420*12 +: 12], 6, 36, SADValues[357*12 +: 12], 5, 37, comp470minVal, comp470minI, comp470minJ);
    wire [11:0] comp471minVal;
    wire [5:0] comp471minI, comp471minJ;
    Comparator comp471(SADValues[294*12 +: 12], 4, 38, SADValues[231*12 +: 12], 3, 39, comp471minVal, comp471minI, comp471minJ);
    wire [11:0] comp472minVal;
    wire [5:0] comp472minI, comp472minJ;
    Comparator comp472(SADValues[168*12 +: 12], 2, 40, SADValues[105*12 +: 12], 1, 41, comp472minVal, comp472minI, comp472minJ);
    wire [11:0] comp473minVal;
    wire [5:0] comp473minI, comp473minJ;
    Comparator comp473(SADValues[42*12 +: 12], 0, 42, SADValues[43*12 +: 12], 0, 43, comp473minVal, comp473minI, comp473minJ);
    wire [11:0] comp474minVal;
    wire [5:0] comp474minI, comp474minJ;
    Comparator comp474(SADValues[106*12 +: 12], 1, 42, SADValues[169*12 +: 12], 2, 41, comp474minVal, comp474minI, comp474minJ);
    wire [11:0] comp475minVal;
    wire [5:0] comp475minI, comp475minJ;
    Comparator comp475(SADValues[232*12 +: 12], 3, 40, SADValues[295*12 +: 12], 4, 39, comp475minVal, comp475minI, comp475minJ);
    wire [11:0] comp476minVal;
    wire [5:0] comp476minI, comp476minJ;
    Comparator comp476(SADValues[358*12 +: 12], 5, 38, SADValues[421*12 +: 12], 6, 37, comp476minVal, comp476minI, comp476minJ);
    wire [11:0] comp477minVal;
    wire [5:0] comp477minI, comp477minJ;
    Comparator comp477(SADValues[484*12 +: 12], 7, 36, SADValues[547*12 +: 12], 8, 35, comp477minVal, comp477minI, comp477minJ);
    wire [11:0] comp478minVal;
    wire [5:0] comp478minI, comp478minJ;
    Comparator comp478(SADValues[610*12 +: 12], 9, 34, SADValues[673*12 +: 12], 10, 33, comp478minVal, comp478minI, comp478minJ);
    wire [11:0] comp479minVal;
    wire [5:0] comp479minI, comp479minJ;
    Comparator comp479(SADValues[736*12 +: 12], 11, 32, SADValues[799*12 +: 12], 12, 31, comp479minVal, comp479minI, comp479minJ);
    wire [11:0] comp480minVal;
    wire [5:0] comp480minI, comp480minJ;
    Comparator comp480(SADValues[862*12 +: 12], 13, 30, SADValues[925*12 +: 12], 14, 29, comp480minVal, comp480minI, comp480minJ);
    wire [11:0] comp481minVal;
    wire [5:0] comp481minI, comp481minJ;
    Comparator comp481(SADValues[988*12 +: 12], 15, 28, SADValues[1051*12 +: 12], 16, 27, comp481minVal, comp481minI, comp481minJ);
    wire [11:0] comp482minVal;
    wire [5:0] comp482minI, comp482minJ;
    Comparator comp482(SADValues[1114*12 +: 12], 17, 26, SADValues[1177*12 +: 12], 18, 25, comp482minVal, comp482minI, comp482minJ);
    wire [11:0] comp483minVal;
    wire [5:0] comp483minI, comp483minJ;
    Comparator comp483(SADValues[1240*12 +: 12], 19, 24, SADValues[1303*12 +: 12], 20, 23, comp483minVal, comp483minI, comp483minJ);
    wire [11:0] comp484minVal;
    wire [5:0] comp484minI, comp484minJ;
    Comparator comp484(SADValues[1366*12 +: 12], 21, 22, SADValues[1429*12 +: 12], 22, 21, comp484minVal, comp484minI, comp484minJ);
    wire [11:0] comp485minVal;
    wire [5:0] comp485minI, comp485minJ;
    Comparator comp485(SADValues[1492*12 +: 12], 23, 20, SADValues[1555*12 +: 12], 24, 19, comp485minVal, comp485minI, comp485minJ);
    wire [11:0] comp486minVal;
    wire [5:0] comp486minI, comp486minJ;
    Comparator comp486(SADValues[1618*12 +: 12], 25, 18, SADValues[1681*12 +: 12], 26, 17, comp486minVal, comp486minI, comp486minJ);
    wire [11:0] comp487minVal;
    wire [5:0] comp487minI, comp487minJ;
    Comparator comp487(SADValues[1744*12 +: 12], 27, 16, SADValues[1807*12 +: 12], 28, 15, comp487minVal, comp487minI, comp487minJ);
    wire [11:0] comp488minVal;
    wire [5:0] comp488minI, comp488minJ;
    Comparator comp488(SADValues[1870*12 +: 12], 29, 14, SADValues[1933*12 +: 12], 30, 13, comp488minVal, comp488minI, comp488minJ);
    wire [11:0] comp489minVal;
    wire [5:0] comp489minI, comp489minJ;
    Comparator comp489(SADValues[1996*12 +: 12], 31, 12, SADValues[2059*12 +: 12], 32, 11, comp489minVal, comp489minI, comp489minJ);
    wire [11:0] comp490minVal;
    wire [5:0] comp490minI, comp490minJ;
    Comparator comp490(SADValues[2122*12 +: 12], 33, 10, SADValues[2185*12 +: 12], 34, 9, comp490minVal, comp490minI, comp490minJ);
    wire [11:0] comp491minVal;
    wire [5:0] comp491minI, comp491minJ;
    Comparator comp491(SADValues[2248*12 +: 12], 35, 8, SADValues[2311*12 +: 12], 36, 7, comp491minVal, comp491minI, comp491minJ);
    wire [11:0] comp492minVal;
    wire [5:0] comp492minI, comp492minJ;
    Comparator comp492(SADValues[2374*12 +: 12], 37, 6, SADValues[2437*12 +: 12], 38, 5, comp492minVal, comp492minI, comp492minJ);
    wire [11:0] comp493minVal;
    wire [5:0] comp493minI, comp493minJ;
    Comparator comp493(SADValues[2500*12 +: 12], 39, 4, SADValues[2563*12 +: 12], 40, 3, comp493minVal, comp493minI, comp493minJ);
    wire [11:0] comp494minVal;
    wire [5:0] comp494minI, comp494minJ;
    Comparator comp494(SADValues[2626*12 +: 12], 41, 2, SADValues[2689*12 +: 12], 42, 1, comp494minVal, comp494minI, comp494minJ);
    wire [11:0] comp495minVal;
    wire [5:0] comp495minI, comp495minJ;
    Comparator comp495(SADValues[2752*12 +: 12], 43, 0, SADValues[2816*12 +: 12], 44, 0, comp495minVal, comp495minI, comp495minJ);
    wire [11:0] comp496minVal;
    wire [5:0] comp496minI, comp496minJ;
    Comparator comp496(SADValues[2753*12 +: 12], 43, 1, SADValues[2690*12 +: 12], 42, 2, comp496minVal, comp496minI, comp496minJ);
    wire [11:0] comp497minVal;
    wire [5:0] comp497minI, comp497minJ;
    Comparator comp497(SADValues[2627*12 +: 12], 41, 3, SADValues[2564*12 +: 12], 40, 4, comp497minVal, comp497minI, comp497minJ);
    wire [11:0] comp498minVal;
    wire [5:0] comp498minI, comp498minJ;
    Comparator comp498(SADValues[2501*12 +: 12], 39, 5, SADValues[2438*12 +: 12], 38, 6, comp498minVal, comp498minI, comp498minJ);
    wire [11:0] comp499minVal;
    wire [5:0] comp499minI, comp499minJ;
    Comparator comp499(SADValues[2375*12 +: 12], 37, 7, SADValues[2312*12 +: 12], 36, 8, comp499minVal, comp499minI, comp499minJ);
    wire [11:0] comp500minVal;
    wire [5:0] comp500minI, comp500minJ;
    Comparator comp500(SADValues[2249*12 +: 12], 35, 9, SADValues[2186*12 +: 12], 34, 10, comp500minVal, comp500minI, comp500minJ);
    wire [11:0] comp501minVal;
    wire [5:0] comp501minI, comp501minJ;
    Comparator comp501(SADValues[2123*12 +: 12], 33, 11, SADValues[2060*12 +: 12], 32, 12, comp501minVal, comp501minI, comp501minJ);
    wire [11:0] comp502minVal;
    wire [5:0] comp502minI, comp502minJ;
    Comparator comp502(SADValues[1997*12 +: 12], 31, 13, SADValues[1934*12 +: 12], 30, 14, comp502minVal, comp502minI, comp502minJ);
    wire [11:0] comp503minVal;
    wire [5:0] comp503minI, comp503minJ;
    Comparator comp503(SADValues[1871*12 +: 12], 29, 15, SADValues[1808*12 +: 12], 28, 16, comp503minVal, comp503minI, comp503minJ);
    wire [11:0] comp504minVal;
    wire [5:0] comp504minI, comp504minJ;
    Comparator comp504(SADValues[1745*12 +: 12], 27, 17, SADValues[1682*12 +: 12], 26, 18, comp504minVal, comp504minI, comp504minJ);
    wire [11:0] comp505minVal;
    wire [5:0] comp505minI, comp505minJ;
    Comparator comp505(SADValues[1619*12 +: 12], 25, 19, SADValues[1556*12 +: 12], 24, 20, comp505minVal, comp505minI, comp505minJ);
    wire [11:0] comp506minVal;
    wire [5:0] comp506minI, comp506minJ;
    Comparator comp506(SADValues[1493*12 +: 12], 23, 21, SADValues[1430*12 +: 12], 22, 22, comp506minVal, comp506minI, comp506minJ);
    wire [11:0] comp507minVal;
    wire [5:0] comp507minI, comp507minJ;
    Comparator comp507(SADValues[1367*12 +: 12], 21, 23, SADValues[1304*12 +: 12], 20, 24, comp507minVal, comp507minI, comp507minJ);
    wire [11:0] comp508minVal;
    wire [5:0] comp508minI, comp508minJ;
    Comparator comp508(SADValues[1241*12 +: 12], 19, 25, SADValues[1178*12 +: 12], 18, 26, comp508minVal, comp508minI, comp508minJ);
    wire [11:0] comp509minVal;
    wire [5:0] comp509minI, comp509minJ;
    Comparator comp509(SADValues[1115*12 +: 12], 17, 27, SADValues[1052*12 +: 12], 16, 28, comp509minVal, comp509minI, comp509minJ);
    wire [11:0] comp510minVal;
    wire [5:0] comp510minI, comp510minJ;
    Comparator comp510(SADValues[989*12 +: 12], 15, 29, SADValues[926*12 +: 12], 14, 30, comp510minVal, comp510minI, comp510minJ);
    wire [11:0] comp511minVal;
    wire [5:0] comp511minI, comp511minJ;
    Comparator comp511(SADValues[863*12 +: 12], 13, 31, SADValues[800*12 +: 12], 12, 32, comp511minVal, comp511minI, comp511minJ);
    wire [11:0] comp512minVal;
    wire [5:0] comp512minI, comp512minJ;
    Comparator comp512(SADValues[737*12 +: 12], 11, 33, SADValues[674*12 +: 12], 10, 34, comp512minVal, comp512minI, comp512minJ);
    wire [11:0] comp513minVal;
    wire [5:0] comp513minI, comp513minJ;
    Comparator comp513(SADValues[611*12 +: 12], 9, 35, SADValues[548*12 +: 12], 8, 36, comp513minVal, comp513minI, comp513minJ);
    wire [11:0] comp514minVal;
    wire [5:0] comp514minI, comp514minJ;
    Comparator comp514(SADValues[485*12 +: 12], 7, 37, SADValues[422*12 +: 12], 6, 38, comp514minVal, comp514minI, comp514minJ);
    wire [11:0] comp515minVal;
    wire [5:0] comp515minI, comp515minJ;
    Comparator comp515(SADValues[359*12 +: 12], 5, 39, SADValues[296*12 +: 12], 4, 40, comp515minVal, comp515minI, comp515minJ);
    wire [11:0] comp516minVal;
    wire [5:0] comp516minI, comp516minJ;
    Comparator comp516(SADValues[233*12 +: 12], 3, 41, SADValues[170*12 +: 12], 2, 42, comp516minVal, comp516minI, comp516minJ);
    wire [11:0] comp517minVal;
    wire [5:0] comp517minI, comp517minJ;
    Comparator comp517(SADValues[107*12 +: 12], 1, 43, SADValues[44*12 +: 12], 0, 44, comp517minVal, comp517minI, comp517minJ);
    wire [11:0] comp518minVal;
    wire [5:0] comp518minI, comp518minJ;
    Comparator comp518(SADValues[45*12 +: 12], 0, 45, SADValues[108*12 +: 12], 1, 44, comp518minVal, comp518minI, comp518minJ);
    wire [11:0] comp519minVal;
    wire [5:0] comp519minI, comp519minJ;
    Comparator comp519(SADValues[171*12 +: 12], 2, 43, SADValues[234*12 +: 12], 3, 42, comp519minVal, comp519minI, comp519minJ);
    wire [11:0] comp520minVal;
    wire [5:0] comp520minI, comp520minJ;
    Comparator comp520(SADValues[297*12 +: 12], 4, 41, SADValues[360*12 +: 12], 5, 40, comp520minVal, comp520minI, comp520minJ);
    wire [11:0] comp521minVal;
    wire [5:0] comp521minI, comp521minJ;
    Comparator comp521(SADValues[423*12 +: 12], 6, 39, SADValues[486*12 +: 12], 7, 38, comp521minVal, comp521minI, comp521minJ);
    wire [11:0] comp522minVal;
    wire [5:0] comp522minI, comp522minJ;
    Comparator comp522(SADValues[549*12 +: 12], 8, 37, SADValues[612*12 +: 12], 9, 36, comp522minVal, comp522minI, comp522minJ);
    wire [11:0] comp523minVal;
    wire [5:0] comp523minI, comp523minJ;
    Comparator comp523(SADValues[675*12 +: 12], 10, 35, SADValues[738*12 +: 12], 11, 34, comp523minVal, comp523minI, comp523minJ);
    wire [11:0] comp524minVal;
    wire [5:0] comp524minI, comp524minJ;
    Comparator comp524(SADValues[801*12 +: 12], 12, 33, SADValues[864*12 +: 12], 13, 32, comp524minVal, comp524minI, comp524minJ);
    wire [11:0] comp525minVal;
    wire [5:0] comp525minI, comp525minJ;
    Comparator comp525(SADValues[927*12 +: 12], 14, 31, SADValues[990*12 +: 12], 15, 30, comp525minVal, comp525minI, comp525minJ);
    wire [11:0] comp526minVal;
    wire [5:0] comp526minI, comp526minJ;
    Comparator comp526(SADValues[1053*12 +: 12], 16, 29, SADValues[1116*12 +: 12], 17, 28, comp526minVal, comp526minI, comp526minJ);
    wire [11:0] comp527minVal;
    wire [5:0] comp527minI, comp527minJ;
    Comparator comp527(SADValues[1179*12 +: 12], 18, 27, SADValues[1242*12 +: 12], 19, 26, comp527minVal, comp527minI, comp527minJ);
    wire [11:0] comp528minVal;
    wire [5:0] comp528minI, comp528minJ;
    Comparator comp528(SADValues[1305*12 +: 12], 20, 25, SADValues[1368*12 +: 12], 21, 24, comp528minVal, comp528minI, comp528minJ);
    wire [11:0] comp529minVal;
    wire [5:0] comp529minI, comp529minJ;
    Comparator comp529(SADValues[1431*12 +: 12], 22, 23, SADValues[1494*12 +: 12], 23, 22, comp529minVal, comp529minI, comp529minJ);
    wire [11:0] comp530minVal;
    wire [5:0] comp530minI, comp530minJ;
    Comparator comp530(SADValues[1557*12 +: 12], 24, 21, SADValues[1620*12 +: 12], 25, 20, comp530minVal, comp530minI, comp530minJ);
    wire [11:0] comp531minVal;
    wire [5:0] comp531minI, comp531minJ;
    Comparator comp531(SADValues[1683*12 +: 12], 26, 19, SADValues[1746*12 +: 12], 27, 18, comp531minVal, comp531minI, comp531minJ);
    wire [11:0] comp532minVal;
    wire [5:0] comp532minI, comp532minJ;
    Comparator comp532(SADValues[1809*12 +: 12], 28, 17, SADValues[1872*12 +: 12], 29, 16, comp532minVal, comp532minI, comp532minJ);
    wire [11:0] comp533minVal;
    wire [5:0] comp533minI, comp533minJ;
    Comparator comp533(SADValues[1935*12 +: 12], 30, 15, SADValues[1998*12 +: 12], 31, 14, comp533minVal, comp533minI, comp533minJ);
    wire [11:0] comp534minVal;
    wire [5:0] comp534minI, comp534minJ;
    Comparator comp534(SADValues[2061*12 +: 12], 32, 13, SADValues[2124*12 +: 12], 33, 12, comp534minVal, comp534minI, comp534minJ);
    wire [11:0] comp535minVal;
    wire [5:0] comp535minI, comp535minJ;
    Comparator comp535(SADValues[2187*12 +: 12], 34, 11, SADValues[2250*12 +: 12], 35, 10, comp535minVal, comp535minI, comp535minJ);
    wire [11:0] comp536minVal;
    wire [5:0] comp536minI, comp536minJ;
    Comparator comp536(SADValues[2313*12 +: 12], 36, 9, SADValues[2376*12 +: 12], 37, 8, comp536minVal, comp536minI, comp536minJ);
    wire [11:0] comp537minVal;
    wire [5:0] comp537minI, comp537minJ;
    Comparator comp537(SADValues[2439*12 +: 12], 38, 7, SADValues[2502*12 +: 12], 39, 6, comp537minVal, comp537minI, comp537minJ);
    wire [11:0] comp538minVal;
    wire [5:0] comp538minI, comp538minJ;
    Comparator comp538(SADValues[2565*12 +: 12], 40, 5, SADValues[2628*12 +: 12], 41, 4, comp538minVal, comp538minI, comp538minJ);
    wire [11:0] comp539minVal;
    wire [5:0] comp539minI, comp539minJ;
    Comparator comp539(SADValues[2691*12 +: 12], 42, 3, SADValues[2754*12 +: 12], 43, 2, comp539minVal, comp539minI, comp539minJ);
    wire [11:0] comp540minVal;
    wire [5:0] comp540minI, comp540minJ;
    Comparator comp540(SADValues[2817*12 +: 12], 44, 1, SADValues[2880*12 +: 12], 45, 0, comp540minVal, comp540minI, comp540minJ);
    wire [11:0] comp541minVal;
    wire [5:0] comp541minI, comp541minJ;
    Comparator comp541(SADValues[2944*12 +: 12], 46, 0, SADValues[2881*12 +: 12], 45, 1, comp541minVal, comp541minI, comp541minJ);
    wire [11:0] comp542minVal;
    wire [5:0] comp542minI, comp542minJ;
    Comparator comp542(SADValues[2818*12 +: 12], 44, 2, SADValues[2755*12 +: 12], 43, 3, comp542minVal, comp542minI, comp542minJ);
    wire [11:0] comp543minVal;
    wire [5:0] comp543minI, comp543minJ;
    Comparator comp543(SADValues[2692*12 +: 12], 42, 4, SADValues[2629*12 +: 12], 41, 5, comp543minVal, comp543minI, comp543minJ);
    wire [11:0] comp544minVal;
    wire [5:0] comp544minI, comp544minJ;
    Comparator comp544(SADValues[2566*12 +: 12], 40, 6, SADValues[2503*12 +: 12], 39, 7, comp544minVal, comp544minI, comp544minJ);
    wire [11:0] comp545minVal;
    wire [5:0] comp545minI, comp545minJ;
    Comparator comp545(SADValues[2440*12 +: 12], 38, 8, SADValues[2377*12 +: 12], 37, 9, comp545minVal, comp545minI, comp545minJ);
    wire [11:0] comp546minVal;
    wire [5:0] comp546minI, comp546minJ;
    Comparator comp546(SADValues[2314*12 +: 12], 36, 10, SADValues[2251*12 +: 12], 35, 11, comp546minVal, comp546minI, comp546minJ);
    wire [11:0] comp547minVal;
    wire [5:0] comp547minI, comp547minJ;
    Comparator comp547(SADValues[2188*12 +: 12], 34, 12, SADValues[2125*12 +: 12], 33, 13, comp547minVal, comp547minI, comp547minJ);
    wire [11:0] comp548minVal;
    wire [5:0] comp548minI, comp548minJ;
    Comparator comp548(SADValues[2062*12 +: 12], 32, 14, SADValues[1999*12 +: 12], 31, 15, comp548minVal, comp548minI, comp548minJ);
    wire [11:0] comp549minVal;
    wire [5:0] comp549minI, comp549minJ;
    Comparator comp549(SADValues[1936*12 +: 12], 30, 16, SADValues[1873*12 +: 12], 29, 17, comp549minVal, comp549minI, comp549minJ);
    wire [11:0] comp550minVal;
    wire [5:0] comp550minI, comp550minJ;
    Comparator comp550(SADValues[1810*12 +: 12], 28, 18, SADValues[1747*12 +: 12], 27, 19, comp550minVal, comp550minI, comp550minJ);
    wire [11:0] comp551minVal;
    wire [5:0] comp551minI, comp551minJ;
    Comparator comp551(SADValues[1684*12 +: 12], 26, 20, SADValues[1621*12 +: 12], 25, 21, comp551minVal, comp551minI, comp551minJ);
    wire [11:0] comp552minVal;
    wire [5:0] comp552minI, comp552minJ;
    Comparator comp552(SADValues[1558*12 +: 12], 24, 22, SADValues[1495*12 +: 12], 23, 23, comp552minVal, comp552minI, comp552minJ);
    wire [11:0] comp553minVal;
    wire [5:0] comp553minI, comp553minJ;
    Comparator comp553(SADValues[1432*12 +: 12], 22, 24, SADValues[1369*12 +: 12], 21, 25, comp553minVal, comp553minI, comp553minJ);
    wire [11:0] comp554minVal;
    wire [5:0] comp554minI, comp554minJ;
    Comparator comp554(SADValues[1306*12 +: 12], 20, 26, SADValues[1243*12 +: 12], 19, 27, comp554minVal, comp554minI, comp554minJ);
    wire [11:0] comp555minVal;
    wire [5:0] comp555minI, comp555minJ;
    Comparator comp555(SADValues[1180*12 +: 12], 18, 28, SADValues[1117*12 +: 12], 17, 29, comp555minVal, comp555minI, comp555minJ);
    wire [11:0] comp556minVal;
    wire [5:0] comp556minI, comp556minJ;
    Comparator comp556(SADValues[1054*12 +: 12], 16, 30, SADValues[991*12 +: 12], 15, 31, comp556minVal, comp556minI, comp556minJ);
    wire [11:0] comp557minVal;
    wire [5:0] comp557minI, comp557minJ;
    Comparator comp557(SADValues[928*12 +: 12], 14, 32, SADValues[865*12 +: 12], 13, 33, comp557minVal, comp557minI, comp557minJ);
    wire [11:0] comp558minVal;
    wire [5:0] comp558minI, comp558minJ;
    Comparator comp558(SADValues[802*12 +: 12], 12, 34, SADValues[739*12 +: 12], 11, 35, comp558minVal, comp558minI, comp558minJ);
    wire [11:0] comp559minVal;
    wire [5:0] comp559minI, comp559minJ;
    Comparator comp559(SADValues[676*12 +: 12], 10, 36, SADValues[613*12 +: 12], 9, 37, comp559minVal, comp559minI, comp559minJ);
    wire [11:0] comp560minVal;
    wire [5:0] comp560minI, comp560minJ;
    Comparator comp560(SADValues[550*12 +: 12], 8, 38, SADValues[487*12 +: 12], 7, 39, comp560minVal, comp560minI, comp560minJ);
    wire [11:0] comp561minVal;
    wire [5:0] comp561minI, comp561minJ;
    Comparator comp561(SADValues[424*12 +: 12], 6, 40, SADValues[361*12 +: 12], 5, 41, comp561minVal, comp561minI, comp561minJ);
    wire [11:0] comp562minVal;
    wire [5:0] comp562minI, comp562minJ;
    Comparator comp562(SADValues[298*12 +: 12], 4, 42, SADValues[235*12 +: 12], 3, 43, comp562minVal, comp562minI, comp562minJ);
    wire [11:0] comp563minVal;
    wire [5:0] comp563minI, comp563minJ;
    Comparator comp563(SADValues[172*12 +: 12], 2, 44, SADValues[109*12 +: 12], 1, 45, comp563minVal, comp563minI, comp563minJ);
    wire [11:0] comp564minVal;
    wire [5:0] comp564minI, comp564minJ;
    Comparator comp564(SADValues[46*12 +: 12], 0, 46, SADValues[47*12 +: 12], 0, 47, comp564minVal, comp564minI, comp564minJ);
    wire [11:0] comp565minVal;
    wire [5:0] comp565minI, comp565minJ;
    Comparator comp565(SADValues[110*12 +: 12], 1, 46, SADValues[173*12 +: 12], 2, 45, comp565minVal, comp565minI, comp565minJ);
    wire [11:0] comp566minVal;
    wire [5:0] comp566minI, comp566minJ;
    Comparator comp566(SADValues[236*12 +: 12], 3, 44, SADValues[299*12 +: 12], 4, 43, comp566minVal, comp566minI, comp566minJ);
    wire [11:0] comp567minVal;
    wire [5:0] comp567minI, comp567minJ;
    Comparator comp567(SADValues[362*12 +: 12], 5, 42, SADValues[425*12 +: 12], 6, 41, comp567minVal, comp567minI, comp567minJ);
    wire [11:0] comp568minVal;
    wire [5:0] comp568minI, comp568minJ;
    Comparator comp568(SADValues[488*12 +: 12], 7, 40, SADValues[551*12 +: 12], 8, 39, comp568minVal, comp568minI, comp568minJ);
    wire [11:0] comp569minVal;
    wire [5:0] comp569minI, comp569minJ;
    Comparator comp569(SADValues[614*12 +: 12], 9, 38, SADValues[677*12 +: 12], 10, 37, comp569minVal, comp569minI, comp569minJ);
    wire [11:0] comp570minVal;
    wire [5:0] comp570minI, comp570minJ;
    Comparator comp570(SADValues[740*12 +: 12], 11, 36, SADValues[803*12 +: 12], 12, 35, comp570minVal, comp570minI, comp570minJ);
    wire [11:0] comp571minVal;
    wire [5:0] comp571minI, comp571minJ;
    Comparator comp571(SADValues[866*12 +: 12], 13, 34, SADValues[929*12 +: 12], 14, 33, comp571minVal, comp571minI, comp571minJ);
    wire [11:0] comp572minVal;
    wire [5:0] comp572minI, comp572minJ;
    Comparator comp572(SADValues[992*12 +: 12], 15, 32, SADValues[1055*12 +: 12], 16, 31, comp572minVal, comp572minI, comp572minJ);
    wire [11:0] comp573minVal;
    wire [5:0] comp573minI, comp573minJ;
    Comparator comp573(SADValues[1118*12 +: 12], 17, 30, SADValues[1181*12 +: 12], 18, 29, comp573minVal, comp573minI, comp573minJ);
    wire [11:0] comp574minVal;
    wire [5:0] comp574minI, comp574minJ;
    Comparator comp574(SADValues[1244*12 +: 12], 19, 28, SADValues[1307*12 +: 12], 20, 27, comp574minVal, comp574minI, comp574minJ);
    wire [11:0] comp575minVal;
    wire [5:0] comp575minI, comp575minJ;
    Comparator comp575(SADValues[1370*12 +: 12], 21, 26, SADValues[1433*12 +: 12], 22, 25, comp575minVal, comp575minI, comp575minJ);
    wire [11:0] comp576minVal;
    wire [5:0] comp576minI, comp576minJ;
    Comparator comp576(SADValues[1496*12 +: 12], 23, 24, SADValues[1559*12 +: 12], 24, 23, comp576minVal, comp576minI, comp576minJ);
    wire [11:0] comp577minVal;
    wire [5:0] comp577minI, comp577minJ;
    Comparator comp577(SADValues[1622*12 +: 12], 25, 22, SADValues[1685*12 +: 12], 26, 21, comp577minVal, comp577minI, comp577minJ);
    wire [11:0] comp578minVal;
    wire [5:0] comp578minI, comp578minJ;
    Comparator comp578(SADValues[1748*12 +: 12], 27, 20, SADValues[1811*12 +: 12], 28, 19, comp578minVal, comp578minI, comp578minJ);
    wire [11:0] comp579minVal;
    wire [5:0] comp579minI, comp579minJ;
    Comparator comp579(SADValues[1874*12 +: 12], 29, 18, SADValues[1937*12 +: 12], 30, 17, comp579minVal, comp579minI, comp579minJ);
    wire [11:0] comp580minVal;
    wire [5:0] comp580minI, comp580minJ;
    Comparator comp580(SADValues[2000*12 +: 12], 31, 16, SADValues[2063*12 +: 12], 32, 15, comp580minVal, comp580minI, comp580minJ);
    wire [11:0] comp581minVal;
    wire [5:0] comp581minI, comp581minJ;
    Comparator comp581(SADValues[2126*12 +: 12], 33, 14, SADValues[2189*12 +: 12], 34, 13, comp581minVal, comp581minI, comp581minJ);
    wire [11:0] comp582minVal;
    wire [5:0] comp582minI, comp582minJ;
    Comparator comp582(SADValues[2252*12 +: 12], 35, 12, SADValues[2315*12 +: 12], 36, 11, comp582minVal, comp582minI, comp582minJ);
    wire [11:0] comp583minVal;
    wire [5:0] comp583minI, comp583minJ;
    Comparator comp583(SADValues[2378*12 +: 12], 37, 10, SADValues[2441*12 +: 12], 38, 9, comp583minVal, comp583minI, comp583minJ);
    wire [11:0] comp584minVal;
    wire [5:0] comp584minI, comp584minJ;
    Comparator comp584(SADValues[2504*12 +: 12], 39, 8, SADValues[2567*12 +: 12], 40, 7, comp584minVal, comp584minI, comp584minJ);
    wire [11:0] comp585minVal;
    wire [5:0] comp585minI, comp585minJ;
    Comparator comp585(SADValues[2630*12 +: 12], 41, 6, SADValues[2693*12 +: 12], 42, 5, comp585minVal, comp585minI, comp585minJ);
    wire [11:0] comp586minVal;
    wire [5:0] comp586minI, comp586minJ;
    Comparator comp586(SADValues[2756*12 +: 12], 43, 4, SADValues[2819*12 +: 12], 44, 3, comp586minVal, comp586minI, comp586minJ);
    wire [11:0] comp587minVal;
    wire [5:0] comp587minI, comp587minJ;
    Comparator comp587(SADValues[2882*12 +: 12], 45, 2, SADValues[2945*12 +: 12], 46, 1, comp587minVal, comp587minI, comp587minJ);
    wire [11:0] comp588minVal;
    wire [5:0] comp588minI, comp588minJ;
    Comparator comp588(SADValues[3008*12 +: 12], 47, 0, SADValues[3072*12 +: 12], 48, 0, comp588minVal, comp588minI, comp588minJ);
    wire [11:0] comp589minVal;
    wire [5:0] comp589minI, comp589minJ;
    Comparator comp589(SADValues[3009*12 +: 12], 47, 1, SADValues[2946*12 +: 12], 46, 2, comp589minVal, comp589minI, comp589minJ);
    wire [11:0] comp590minVal;
    wire [5:0] comp590minI, comp590minJ;
    Comparator comp590(SADValues[2883*12 +: 12], 45, 3, SADValues[2820*12 +: 12], 44, 4, comp590minVal, comp590minI, comp590minJ);
    wire [11:0] comp591minVal;
    wire [5:0] comp591minI, comp591minJ;
    Comparator comp591(SADValues[2757*12 +: 12], 43, 5, SADValues[2694*12 +: 12], 42, 6, comp591minVal, comp591minI, comp591minJ);
    wire [11:0] comp592minVal;
    wire [5:0] comp592minI, comp592minJ;
    Comparator comp592(SADValues[2631*12 +: 12], 41, 7, SADValues[2568*12 +: 12], 40, 8, comp592minVal, comp592minI, comp592minJ);
    wire [11:0] comp593minVal;
    wire [5:0] comp593minI, comp593minJ;
    Comparator comp593(SADValues[2505*12 +: 12], 39, 9, SADValues[2442*12 +: 12], 38, 10, comp593minVal, comp593minI, comp593minJ);
    wire [11:0] comp594minVal;
    wire [5:0] comp594minI, comp594minJ;
    Comparator comp594(SADValues[2379*12 +: 12], 37, 11, SADValues[2316*12 +: 12], 36, 12, comp594minVal, comp594minI, comp594minJ);
    wire [11:0] comp595minVal;
    wire [5:0] comp595minI, comp595minJ;
    Comparator comp595(SADValues[2253*12 +: 12], 35, 13, SADValues[2190*12 +: 12], 34, 14, comp595minVal, comp595minI, comp595minJ);
    wire [11:0] comp596minVal;
    wire [5:0] comp596minI, comp596minJ;
    Comparator comp596(SADValues[2127*12 +: 12], 33, 15, SADValues[2064*12 +: 12], 32, 16, comp596minVal, comp596minI, comp596minJ);
    wire [11:0] comp597minVal;
    wire [5:0] comp597minI, comp597minJ;
    Comparator comp597(SADValues[2001*12 +: 12], 31, 17, SADValues[1938*12 +: 12], 30, 18, comp597minVal, comp597minI, comp597minJ);
    wire [11:0] comp598minVal;
    wire [5:0] comp598minI, comp598minJ;
    Comparator comp598(SADValues[1875*12 +: 12], 29, 19, SADValues[1812*12 +: 12], 28, 20, comp598minVal, comp598minI, comp598minJ);
    wire [11:0] comp599minVal;
    wire [5:0] comp599minI, comp599minJ;
    Comparator comp599(SADValues[1749*12 +: 12], 27, 21, SADValues[1686*12 +: 12], 26, 22, comp599minVal, comp599minI, comp599minJ);
    wire [11:0] comp600minVal;
    wire [5:0] comp600minI, comp600minJ;
    Comparator comp600(SADValues[1623*12 +: 12], 25, 23, SADValues[1560*12 +: 12], 24, 24, comp600minVal, comp600minI, comp600minJ);
    wire [11:0] comp601minVal;
    wire [5:0] comp601minI, comp601minJ;
    Comparator comp601(SADValues[1497*12 +: 12], 23, 25, SADValues[1434*12 +: 12], 22, 26, comp601minVal, comp601minI, comp601minJ);
    wire [11:0] comp602minVal;
    wire [5:0] comp602minI, comp602minJ;
    Comparator comp602(SADValues[1371*12 +: 12], 21, 27, SADValues[1308*12 +: 12], 20, 28, comp602minVal, comp602minI, comp602minJ);
    wire [11:0] comp603minVal;
    wire [5:0] comp603minI, comp603minJ;
    Comparator comp603(SADValues[1245*12 +: 12], 19, 29, SADValues[1182*12 +: 12], 18, 30, comp603minVal, comp603minI, comp603minJ);
    wire [11:0] comp604minVal;
    wire [5:0] comp604minI, comp604minJ;
    Comparator comp604(SADValues[1119*12 +: 12], 17, 31, SADValues[1056*12 +: 12], 16, 32, comp604minVal, comp604minI, comp604minJ);
    wire [11:0] comp605minVal;
    wire [5:0] comp605minI, comp605minJ;
    Comparator comp605(SADValues[993*12 +: 12], 15, 33, SADValues[930*12 +: 12], 14, 34, comp605minVal, comp605minI, comp605minJ);
    wire [11:0] comp606minVal;
    wire [5:0] comp606minI, comp606minJ;
    Comparator comp606(SADValues[867*12 +: 12], 13, 35, SADValues[804*12 +: 12], 12, 36, comp606minVal, comp606minI, comp606minJ);
    wire [11:0] comp607minVal;
    wire [5:0] comp607minI, comp607minJ;
    Comparator comp607(SADValues[741*12 +: 12], 11, 37, SADValues[678*12 +: 12], 10, 38, comp607minVal, comp607minI, comp607minJ);
    wire [11:0] comp608minVal;
    wire [5:0] comp608minI, comp608minJ;
    Comparator comp608(SADValues[615*12 +: 12], 9, 39, SADValues[552*12 +: 12], 8, 40, comp608minVal, comp608minI, comp608minJ);
    wire [11:0] comp609minVal;
    wire [5:0] comp609minI, comp609minJ;
    Comparator comp609(SADValues[489*12 +: 12], 7, 41, SADValues[426*12 +: 12], 6, 42, comp609minVal, comp609minI, comp609minJ);
    wire [11:0] comp610minVal;
    wire [5:0] comp610minI, comp610minJ;
    Comparator comp610(SADValues[363*12 +: 12], 5, 43, SADValues[300*12 +: 12], 4, 44, comp610minVal, comp610minI, comp610minJ);
    wire [11:0] comp611minVal;
    wire [5:0] comp611minI, comp611minJ;
    Comparator comp611(SADValues[237*12 +: 12], 3, 45, SADValues[174*12 +: 12], 2, 46, comp611minVal, comp611minI, comp611minJ);
    wire [11:0] comp612minVal;
    wire [5:0] comp612minI, comp612minJ;
    Comparator comp612(SADValues[111*12 +: 12], 1, 47, SADValues[48*12 +: 12], 0, 48, comp612minVal, comp612minI, comp612minJ);
    wire [11:0] comp613minVal;
    wire [5:0] comp613minI, comp613minJ;
    Comparator comp613(SADValues[49*12 +: 12], 0, 49, SADValues[112*12 +: 12], 1, 48, comp613minVal, comp613minI, comp613minJ);
    wire [11:0] comp614minVal;
    wire [5:0] comp614minI, comp614minJ;
    Comparator comp614(SADValues[175*12 +: 12], 2, 47, SADValues[238*12 +: 12], 3, 46, comp614minVal, comp614minI, comp614minJ);
    wire [11:0] comp615minVal;
    wire [5:0] comp615minI, comp615minJ;
    Comparator comp615(SADValues[301*12 +: 12], 4, 45, SADValues[364*12 +: 12], 5, 44, comp615minVal, comp615minI, comp615minJ);
    wire [11:0] comp616minVal;
    wire [5:0] comp616minI, comp616minJ;
    Comparator comp616(SADValues[427*12 +: 12], 6, 43, SADValues[490*12 +: 12], 7, 42, comp616minVal, comp616minI, comp616minJ);
    wire [11:0] comp617minVal;
    wire [5:0] comp617minI, comp617minJ;
    Comparator comp617(SADValues[553*12 +: 12], 8, 41, SADValues[616*12 +: 12], 9, 40, comp617minVal, comp617minI, comp617minJ);
    wire [11:0] comp618minVal;
    wire [5:0] comp618minI, comp618minJ;
    Comparator comp618(SADValues[679*12 +: 12], 10, 39, SADValues[742*12 +: 12], 11, 38, comp618minVal, comp618minI, comp618minJ);
    wire [11:0] comp619minVal;
    wire [5:0] comp619minI, comp619minJ;
    Comparator comp619(SADValues[805*12 +: 12], 12, 37, SADValues[868*12 +: 12], 13, 36, comp619minVal, comp619minI, comp619minJ);
    wire [11:0] comp620minVal;
    wire [5:0] comp620minI, comp620minJ;
    Comparator comp620(SADValues[931*12 +: 12], 14, 35, SADValues[994*12 +: 12], 15, 34, comp620minVal, comp620minI, comp620minJ);
    wire [11:0] comp621minVal;
    wire [5:0] comp621minI, comp621minJ;
    Comparator comp621(SADValues[1057*12 +: 12], 16, 33, SADValues[1120*12 +: 12], 17, 32, comp621minVal, comp621minI, comp621minJ);
    wire [11:0] comp622minVal;
    wire [5:0] comp622minI, comp622minJ;
    Comparator comp622(SADValues[1183*12 +: 12], 18, 31, SADValues[1246*12 +: 12], 19, 30, comp622minVal, comp622minI, comp622minJ);
    wire [11:0] comp623minVal;
    wire [5:0] comp623minI, comp623minJ;
    Comparator comp623(SADValues[1309*12 +: 12], 20, 29, SADValues[1372*12 +: 12], 21, 28, comp623minVal, comp623minI, comp623minJ);
    wire [11:0] comp624minVal;
    wire [5:0] comp624minI, comp624minJ;
    Comparator comp624(SADValues[1435*12 +: 12], 22, 27, SADValues[1498*12 +: 12], 23, 26, comp624minVal, comp624minI, comp624minJ);
    wire [11:0] comp625minVal;
    wire [5:0] comp625minI, comp625minJ;
    Comparator comp625(SADValues[1561*12 +: 12], 24, 25, SADValues[1624*12 +: 12], 25, 24, comp625minVal, comp625minI, comp625minJ);
    wire [11:0] comp626minVal;
    wire [5:0] comp626minI, comp626minJ;
    Comparator comp626(SADValues[1687*12 +: 12], 26, 23, SADValues[1750*12 +: 12], 27, 22, comp626minVal, comp626minI, comp626minJ);
    wire [11:0] comp627minVal;
    wire [5:0] comp627minI, comp627minJ;
    Comparator comp627(SADValues[1813*12 +: 12], 28, 21, SADValues[1876*12 +: 12], 29, 20, comp627minVal, comp627minI, comp627minJ);
    wire [11:0] comp628minVal;
    wire [5:0] comp628minI, comp628minJ;
    Comparator comp628(SADValues[1939*12 +: 12], 30, 19, SADValues[2002*12 +: 12], 31, 18, comp628minVal, comp628minI, comp628minJ);
    wire [11:0] comp629minVal;
    wire [5:0] comp629minI, comp629minJ;
    Comparator comp629(SADValues[2065*12 +: 12], 32, 17, SADValues[2128*12 +: 12], 33, 16, comp629minVal, comp629minI, comp629minJ);
    wire [11:0] comp630minVal;
    wire [5:0] comp630minI, comp630minJ;
    Comparator comp630(SADValues[2191*12 +: 12], 34, 15, SADValues[2254*12 +: 12], 35, 14, comp630minVal, comp630minI, comp630minJ);
    wire [11:0] comp631minVal;
    wire [5:0] comp631minI, comp631minJ;
    Comparator comp631(SADValues[2317*12 +: 12], 36, 13, SADValues[2380*12 +: 12], 37, 12, comp631minVal, comp631minI, comp631minJ);
    wire [11:0] comp632minVal;
    wire [5:0] comp632minI, comp632minJ;
    Comparator comp632(SADValues[2443*12 +: 12], 38, 11, SADValues[2506*12 +: 12], 39, 10, comp632minVal, comp632minI, comp632minJ);
    wire [11:0] comp633minVal;
    wire [5:0] comp633minI, comp633minJ;
    Comparator comp633(SADValues[2569*12 +: 12], 40, 9, SADValues[2632*12 +: 12], 41, 8, comp633minVal, comp633minI, comp633minJ);
    wire [11:0] comp634minVal;
    wire [5:0] comp634minI, comp634minJ;
    Comparator comp634(SADValues[2695*12 +: 12], 42, 7, SADValues[2758*12 +: 12], 43, 6, comp634minVal, comp634minI, comp634minJ);
    wire [11:0] comp635minVal;
    wire [5:0] comp635minI, comp635minJ;
    Comparator comp635(SADValues[2821*12 +: 12], 44, 5, SADValues[2884*12 +: 12], 45, 4, comp635minVal, comp635minI, comp635minJ);
    wire [11:0] comp636minVal;
    wire [5:0] comp636minI, comp636minJ;
    Comparator comp636(SADValues[2947*12 +: 12], 46, 3, SADValues[3010*12 +: 12], 47, 2, comp636minVal, comp636minI, comp636minJ);
    wire [11:0] comp637minVal;
    wire [5:0] comp637minI, comp637minJ;
    Comparator comp637(SADValues[3073*12 +: 12], 48, 1, SADValues[3136*12 +: 12], 49, 0, comp637minVal, comp637minI, comp637minJ);
    wire [11:0] comp638minVal;
    wire [5:0] comp638minI, comp638minJ;
    Comparator comp638(SADValues[3200*12 +: 12], 50, 0, SADValues[3137*12 +: 12], 49, 1, comp638minVal, comp638minI, comp638minJ);
    wire [11:0] comp639minVal;
    wire [5:0] comp639minI, comp639minJ;
    Comparator comp639(SADValues[3074*12 +: 12], 48, 2, SADValues[3011*12 +: 12], 47, 3, comp639minVal, comp639minI, comp639minJ);
    wire [11:0] comp640minVal;
    wire [5:0] comp640minI, comp640minJ;
    Comparator comp640(SADValues[2948*12 +: 12], 46, 4, SADValues[2885*12 +: 12], 45, 5, comp640minVal, comp640minI, comp640minJ);
    wire [11:0] comp641minVal;
    wire [5:0] comp641minI, comp641minJ;
    Comparator comp641(SADValues[2822*12 +: 12], 44, 6, SADValues[2759*12 +: 12], 43, 7, comp641minVal, comp641minI, comp641minJ);
    wire [11:0] comp642minVal;
    wire [5:0] comp642minI, comp642minJ;
    Comparator comp642(SADValues[2696*12 +: 12], 42, 8, SADValues[2633*12 +: 12], 41, 9, comp642minVal, comp642minI, comp642minJ);
    wire [11:0] comp643minVal;
    wire [5:0] comp643minI, comp643minJ;
    Comparator comp643(SADValues[2570*12 +: 12], 40, 10, SADValues[2507*12 +: 12], 39, 11, comp643minVal, comp643minI, comp643minJ);
    wire [11:0] comp644minVal;
    wire [5:0] comp644minI, comp644minJ;
    Comparator comp644(SADValues[2444*12 +: 12], 38, 12, SADValues[2381*12 +: 12], 37, 13, comp644minVal, comp644minI, comp644minJ);
    wire [11:0] comp645minVal;
    wire [5:0] comp645minI, comp645minJ;
    Comparator comp645(SADValues[2318*12 +: 12], 36, 14, SADValues[2255*12 +: 12], 35, 15, comp645minVal, comp645minI, comp645minJ);
    wire [11:0] comp646minVal;
    wire [5:0] comp646minI, comp646minJ;
    Comparator comp646(SADValues[2192*12 +: 12], 34, 16, SADValues[2129*12 +: 12], 33, 17, comp646minVal, comp646minI, comp646minJ);
    wire [11:0] comp647minVal;
    wire [5:0] comp647minI, comp647minJ;
    Comparator comp647(SADValues[2066*12 +: 12], 32, 18, SADValues[2003*12 +: 12], 31, 19, comp647minVal, comp647minI, comp647minJ);
    wire [11:0] comp648minVal;
    wire [5:0] comp648minI, comp648minJ;
    Comparator comp648(SADValues[1940*12 +: 12], 30, 20, SADValues[1877*12 +: 12], 29, 21, comp648minVal, comp648minI, comp648minJ);
    wire [11:0] comp649minVal;
    wire [5:0] comp649minI, comp649minJ;
    Comparator comp649(SADValues[1814*12 +: 12], 28, 22, SADValues[1751*12 +: 12], 27, 23, comp649minVal, comp649minI, comp649minJ);
    wire [11:0] comp650minVal;
    wire [5:0] comp650minI, comp650minJ;
    Comparator comp650(SADValues[1688*12 +: 12], 26, 24, SADValues[1625*12 +: 12], 25, 25, comp650minVal, comp650minI, comp650minJ);
    wire [11:0] comp651minVal;
    wire [5:0] comp651minI, comp651minJ;
    Comparator comp651(SADValues[1562*12 +: 12], 24, 26, SADValues[1499*12 +: 12], 23, 27, comp651minVal, comp651minI, comp651minJ);
    wire [11:0] comp652minVal;
    wire [5:0] comp652minI, comp652minJ;
    Comparator comp652(SADValues[1436*12 +: 12], 22, 28, SADValues[1373*12 +: 12], 21, 29, comp652minVal, comp652minI, comp652minJ);
    wire [11:0] comp653minVal;
    wire [5:0] comp653minI, comp653minJ;
    Comparator comp653(SADValues[1310*12 +: 12], 20, 30, SADValues[1247*12 +: 12], 19, 31, comp653minVal, comp653minI, comp653minJ);
    wire [11:0] comp654minVal;
    wire [5:0] comp654minI, comp654minJ;
    Comparator comp654(SADValues[1184*12 +: 12], 18, 32, SADValues[1121*12 +: 12], 17, 33, comp654minVal, comp654minI, comp654minJ);
    wire [11:0] comp655minVal;
    wire [5:0] comp655minI, comp655minJ;
    Comparator comp655(SADValues[1058*12 +: 12], 16, 34, SADValues[995*12 +: 12], 15, 35, comp655minVal, comp655minI, comp655minJ);
    wire [11:0] comp656minVal;
    wire [5:0] comp656minI, comp656minJ;
    Comparator comp656(SADValues[932*12 +: 12], 14, 36, SADValues[869*12 +: 12], 13, 37, comp656minVal, comp656minI, comp656minJ);
    wire [11:0] comp657minVal;
    wire [5:0] comp657minI, comp657minJ;
    Comparator comp657(SADValues[806*12 +: 12], 12, 38, SADValues[743*12 +: 12], 11, 39, comp657minVal, comp657minI, comp657minJ);
    wire [11:0] comp658minVal;
    wire [5:0] comp658minI, comp658minJ;
    Comparator comp658(SADValues[680*12 +: 12], 10, 40, SADValues[617*12 +: 12], 9, 41, comp658minVal, comp658minI, comp658minJ);
    wire [11:0] comp659minVal;
    wire [5:0] comp659minI, comp659minJ;
    Comparator comp659(SADValues[554*12 +: 12], 8, 42, SADValues[491*12 +: 12], 7, 43, comp659minVal, comp659minI, comp659minJ);
    wire [11:0] comp660minVal;
    wire [5:0] comp660minI, comp660minJ;
    Comparator comp660(SADValues[428*12 +: 12], 6, 44, SADValues[365*12 +: 12], 5, 45, comp660minVal, comp660minI, comp660minJ);
    wire [11:0] comp661minVal;
    wire [5:0] comp661minI, comp661minJ;
    Comparator comp661(SADValues[302*12 +: 12], 4, 46, SADValues[239*12 +: 12], 3, 47, comp661minVal, comp661minI, comp661minJ);
    wire [11:0] comp662minVal;
    wire [5:0] comp662minI, comp662minJ;
    Comparator comp662(SADValues[176*12 +: 12], 2, 48, SADValues[113*12 +: 12], 1, 49, comp662minVal, comp662minI, comp662minJ);
    wire [11:0] comp663minVal;
    wire [5:0] comp663minI, comp663minJ;
    Comparator comp663(SADValues[50*12 +: 12], 0, 50, SADValues[51*12 +: 12], 0, 51, comp663minVal, comp663minI, comp663minJ);
    wire [11:0] comp664minVal;
    wire [5:0] comp664minI, comp664minJ;
    Comparator comp664(SADValues[114*12 +: 12], 1, 50, SADValues[177*12 +: 12], 2, 49, comp664minVal, comp664minI, comp664minJ);
    wire [11:0] comp665minVal;
    wire [5:0] comp665minI, comp665minJ;
    Comparator comp665(SADValues[240*12 +: 12], 3, 48, SADValues[303*12 +: 12], 4, 47, comp665minVal, comp665minI, comp665minJ);
    wire [11:0] comp666minVal;
    wire [5:0] comp666minI, comp666minJ;
    Comparator comp666(SADValues[366*12 +: 12], 5, 46, SADValues[429*12 +: 12], 6, 45, comp666minVal, comp666minI, comp666minJ);
    wire [11:0] comp667minVal;
    wire [5:0] comp667minI, comp667minJ;
    Comparator comp667(SADValues[492*12 +: 12], 7, 44, SADValues[555*12 +: 12], 8, 43, comp667minVal, comp667minI, comp667minJ);
    wire [11:0] comp668minVal;
    wire [5:0] comp668minI, comp668minJ;
    Comparator comp668(SADValues[618*12 +: 12], 9, 42, SADValues[681*12 +: 12], 10, 41, comp668minVal, comp668minI, comp668minJ);
    wire [11:0] comp669minVal;
    wire [5:0] comp669minI, comp669minJ;
    Comparator comp669(SADValues[744*12 +: 12], 11, 40, SADValues[807*12 +: 12], 12, 39, comp669minVal, comp669minI, comp669minJ);
    wire [11:0] comp670minVal;
    wire [5:0] comp670minI, comp670minJ;
    Comparator comp670(SADValues[870*12 +: 12], 13, 38, SADValues[933*12 +: 12], 14, 37, comp670minVal, comp670minI, comp670minJ);
    wire [11:0] comp671minVal;
    wire [5:0] comp671minI, comp671minJ;
    Comparator comp671(SADValues[996*12 +: 12], 15, 36, SADValues[1059*12 +: 12], 16, 35, comp671minVal, comp671minI, comp671minJ);
    wire [11:0] comp672minVal;
    wire [5:0] comp672minI, comp672minJ;
    Comparator comp672(SADValues[1122*12 +: 12], 17, 34, SADValues[1185*12 +: 12], 18, 33, comp672minVal, comp672minI, comp672minJ);
    wire [11:0] comp673minVal;
    wire [5:0] comp673minI, comp673minJ;
    Comparator comp673(SADValues[1248*12 +: 12], 19, 32, SADValues[1311*12 +: 12], 20, 31, comp673minVal, comp673minI, comp673minJ);
    wire [11:0] comp674minVal;
    wire [5:0] comp674minI, comp674minJ;
    Comparator comp674(SADValues[1374*12 +: 12], 21, 30, SADValues[1437*12 +: 12], 22, 29, comp674minVal, comp674minI, comp674minJ);
    wire [11:0] comp675minVal;
    wire [5:0] comp675minI, comp675minJ;
    Comparator comp675(SADValues[1500*12 +: 12], 23, 28, SADValues[1563*12 +: 12], 24, 27, comp675minVal, comp675minI, comp675minJ);
    wire [11:0] comp676minVal;
    wire [5:0] comp676minI, comp676minJ;
    Comparator comp676(SADValues[1626*12 +: 12], 25, 26, SADValues[1689*12 +: 12], 26, 25, comp676minVal, comp676minI, comp676minJ);
    wire [11:0] comp677minVal;
    wire [5:0] comp677minI, comp677minJ;
    Comparator comp677(SADValues[1752*12 +: 12], 27, 24, SADValues[1815*12 +: 12], 28, 23, comp677minVal, comp677minI, comp677minJ);
    wire [11:0] comp678minVal;
    wire [5:0] comp678minI, comp678minJ;
    Comparator comp678(SADValues[1878*12 +: 12], 29, 22, SADValues[1941*12 +: 12], 30, 21, comp678minVal, comp678minI, comp678minJ);
    wire [11:0] comp679minVal;
    wire [5:0] comp679minI, comp679minJ;
    Comparator comp679(SADValues[2004*12 +: 12], 31, 20, SADValues[2067*12 +: 12], 32, 19, comp679minVal, comp679minI, comp679minJ);
    wire [11:0] comp680minVal;
    wire [5:0] comp680minI, comp680minJ;
    Comparator comp680(SADValues[2130*12 +: 12], 33, 18, SADValues[2193*12 +: 12], 34, 17, comp680minVal, comp680minI, comp680minJ);
    wire [11:0] comp681minVal;
    wire [5:0] comp681minI, comp681minJ;
    Comparator comp681(SADValues[2256*12 +: 12], 35, 16, SADValues[2319*12 +: 12], 36, 15, comp681minVal, comp681minI, comp681minJ);
    wire [11:0] comp682minVal;
    wire [5:0] comp682minI, comp682minJ;
    Comparator comp682(SADValues[2382*12 +: 12], 37, 14, SADValues[2445*12 +: 12], 38, 13, comp682minVal, comp682minI, comp682minJ);
    wire [11:0] comp683minVal;
    wire [5:0] comp683minI, comp683minJ;
    Comparator comp683(SADValues[2508*12 +: 12], 39, 12, SADValues[2571*12 +: 12], 40, 11, comp683minVal, comp683minI, comp683minJ);
    wire [11:0] comp684minVal;
    wire [5:0] comp684minI, comp684minJ;
    Comparator comp684(SADValues[2634*12 +: 12], 41, 10, SADValues[2697*12 +: 12], 42, 9, comp684minVal, comp684minI, comp684minJ);
    wire [11:0] comp685minVal;
    wire [5:0] comp685minI, comp685minJ;
    Comparator comp685(SADValues[2760*12 +: 12], 43, 8, SADValues[2823*12 +: 12], 44, 7, comp685minVal, comp685minI, comp685minJ);
    wire [11:0] comp686minVal;
    wire [5:0] comp686minI, comp686minJ;
    Comparator comp686(SADValues[2886*12 +: 12], 45, 6, SADValues[2949*12 +: 12], 46, 5, comp686minVal, comp686minI, comp686minJ);
    wire [11:0] comp687minVal;
    wire [5:0] comp687minI, comp687minJ;
    Comparator comp687(SADValues[3012*12 +: 12], 47, 4, SADValues[3075*12 +: 12], 48, 3, comp687minVal, comp687minI, comp687minJ);
    wire [11:0] comp688minVal;
    wire [5:0] comp688minI, comp688minJ;
    Comparator comp688(SADValues[3138*12 +: 12], 49, 2, SADValues[3201*12 +: 12], 50, 1, comp688minVal, comp688minI, comp688minJ);
    wire [11:0] comp689minVal;
    wire [5:0] comp689minI, comp689minJ;
    Comparator comp689(SADValues[3264*12 +: 12], 51, 0, SADValues[3328*12 +: 12], 52, 0, comp689minVal, comp689minI, comp689minJ);
    wire [11:0] comp690minVal;
    wire [5:0] comp690minI, comp690minJ;
    Comparator comp690(SADValues[3265*12 +: 12], 51, 1, SADValues[3202*12 +: 12], 50, 2, comp690minVal, comp690minI, comp690minJ);
    wire [11:0] comp691minVal;
    wire [5:0] comp691minI, comp691minJ;
    Comparator comp691(SADValues[3139*12 +: 12], 49, 3, SADValues[3076*12 +: 12], 48, 4, comp691minVal, comp691minI, comp691minJ);
    wire [11:0] comp692minVal;
    wire [5:0] comp692minI, comp692minJ;
    Comparator comp692(SADValues[3013*12 +: 12], 47, 5, SADValues[2950*12 +: 12], 46, 6, comp692minVal, comp692minI, comp692minJ);
    wire [11:0] comp693minVal;
    wire [5:0] comp693minI, comp693minJ;
    Comparator comp693(SADValues[2887*12 +: 12], 45, 7, SADValues[2824*12 +: 12], 44, 8, comp693minVal, comp693minI, comp693minJ);
    wire [11:0] comp694minVal;
    wire [5:0] comp694minI, comp694minJ;
    Comparator comp694(SADValues[2761*12 +: 12], 43, 9, SADValues[2698*12 +: 12], 42, 10, comp694minVal, comp694minI, comp694minJ);
    wire [11:0] comp695minVal;
    wire [5:0] comp695minI, comp695minJ;
    Comparator comp695(SADValues[2635*12 +: 12], 41, 11, SADValues[2572*12 +: 12], 40, 12, comp695minVal, comp695minI, comp695minJ);
    wire [11:0] comp696minVal;
    wire [5:0] comp696minI, comp696minJ;
    Comparator comp696(SADValues[2509*12 +: 12], 39, 13, SADValues[2446*12 +: 12], 38, 14, comp696minVal, comp696minI, comp696minJ);
    wire [11:0] comp697minVal;
    wire [5:0] comp697minI, comp697minJ;
    Comparator comp697(SADValues[2383*12 +: 12], 37, 15, SADValues[2320*12 +: 12], 36, 16, comp697minVal, comp697minI, comp697minJ);
    wire [11:0] comp698minVal;
    wire [5:0] comp698minI, comp698minJ;
    Comparator comp698(SADValues[2257*12 +: 12], 35, 17, SADValues[2194*12 +: 12], 34, 18, comp698minVal, comp698minI, comp698minJ);
    wire [11:0] comp699minVal;
    wire [5:0] comp699minI, comp699minJ;
    Comparator comp699(SADValues[2131*12 +: 12], 33, 19, SADValues[2068*12 +: 12], 32, 20, comp699minVal, comp699minI, comp699minJ);
    wire [11:0] comp700minVal;
    wire [5:0] comp700minI, comp700minJ;
    Comparator comp700(SADValues[2005*12 +: 12], 31, 21, SADValues[1942*12 +: 12], 30, 22, comp700minVal, comp700minI, comp700minJ);
    wire [11:0] comp701minVal;
    wire [5:0] comp701minI, comp701minJ;
    Comparator comp701(SADValues[1879*12 +: 12], 29, 23, SADValues[1816*12 +: 12], 28, 24, comp701minVal, comp701minI, comp701minJ);
    wire [11:0] comp702minVal;
    wire [5:0] comp702minI, comp702minJ;
    Comparator comp702(SADValues[1753*12 +: 12], 27, 25, SADValues[1690*12 +: 12], 26, 26, comp702minVal, comp702minI, comp702minJ);
    wire [11:0] comp703minVal;
    wire [5:0] comp703minI, comp703minJ;
    Comparator comp703(SADValues[1627*12 +: 12], 25, 27, SADValues[1564*12 +: 12], 24, 28, comp703minVal, comp703minI, comp703minJ);
    wire [11:0] comp704minVal;
    wire [5:0] comp704minI, comp704minJ;
    Comparator comp704(SADValues[1501*12 +: 12], 23, 29, SADValues[1438*12 +: 12], 22, 30, comp704minVal, comp704minI, comp704minJ);
    wire [11:0] comp705minVal;
    wire [5:0] comp705minI, comp705minJ;
    Comparator comp705(SADValues[1375*12 +: 12], 21, 31, SADValues[1312*12 +: 12], 20, 32, comp705minVal, comp705minI, comp705minJ);
    wire [11:0] comp706minVal;
    wire [5:0] comp706minI, comp706minJ;
    Comparator comp706(SADValues[1249*12 +: 12], 19, 33, SADValues[1186*12 +: 12], 18, 34, comp706minVal, comp706minI, comp706minJ);
    wire [11:0] comp707minVal;
    wire [5:0] comp707minI, comp707minJ;
    Comparator comp707(SADValues[1123*12 +: 12], 17, 35, SADValues[1060*12 +: 12], 16, 36, comp707minVal, comp707minI, comp707minJ);
    wire [11:0] comp708minVal;
    wire [5:0] comp708minI, comp708minJ;
    Comparator comp708(SADValues[997*12 +: 12], 15, 37, SADValues[934*12 +: 12], 14, 38, comp708minVal, comp708minI, comp708minJ);
    wire [11:0] comp709minVal;
    wire [5:0] comp709minI, comp709minJ;
    Comparator comp709(SADValues[871*12 +: 12], 13, 39, SADValues[808*12 +: 12], 12, 40, comp709minVal, comp709minI, comp709minJ);
    wire [11:0] comp710minVal;
    wire [5:0] comp710minI, comp710minJ;
    Comparator comp710(SADValues[745*12 +: 12], 11, 41, SADValues[682*12 +: 12], 10, 42, comp710minVal, comp710minI, comp710minJ);
    wire [11:0] comp711minVal;
    wire [5:0] comp711minI, comp711minJ;
    Comparator comp711(SADValues[619*12 +: 12], 9, 43, SADValues[556*12 +: 12], 8, 44, comp711minVal, comp711minI, comp711minJ);
    wire [11:0] comp712minVal;
    wire [5:0] comp712minI, comp712minJ;
    Comparator comp712(SADValues[493*12 +: 12], 7, 45, SADValues[430*12 +: 12], 6, 46, comp712minVal, comp712minI, comp712minJ);
    wire [11:0] comp713minVal;
    wire [5:0] comp713minI, comp713minJ;
    Comparator comp713(SADValues[367*12 +: 12], 5, 47, SADValues[304*12 +: 12], 4, 48, comp713minVal, comp713minI, comp713minJ);
    wire [11:0] comp714minVal;
    wire [5:0] comp714minI, comp714minJ;
    Comparator comp714(SADValues[241*12 +: 12], 3, 49, SADValues[178*12 +: 12], 2, 50, comp714minVal, comp714minI, comp714minJ);
    wire [11:0] comp715minVal;
    wire [5:0] comp715minI, comp715minJ;
    Comparator comp715(SADValues[115*12 +: 12], 1, 51, SADValues[52*12 +: 12], 0, 52, comp715minVal, comp715minI, comp715minJ);
    wire [11:0] comp716minVal;
    wire [5:0] comp716minI, comp716minJ;
    Comparator comp716(SADValues[53*12 +: 12], 0, 53, SADValues[116*12 +: 12], 1, 52, comp716minVal, comp716minI, comp716minJ);
    wire [11:0] comp717minVal;
    wire [5:0] comp717minI, comp717minJ;
    Comparator comp717(SADValues[179*12 +: 12], 2, 51, SADValues[242*12 +: 12], 3, 50, comp717minVal, comp717minI, comp717minJ);
    wire [11:0] comp718minVal;
    wire [5:0] comp718minI, comp718minJ;
    Comparator comp718(SADValues[305*12 +: 12], 4, 49, SADValues[368*12 +: 12], 5, 48, comp718minVal, comp718minI, comp718minJ);
    wire [11:0] comp719minVal;
    wire [5:0] comp719minI, comp719minJ;
    Comparator comp719(SADValues[431*12 +: 12], 6, 47, SADValues[494*12 +: 12], 7, 46, comp719minVal, comp719minI, comp719minJ);
    wire [11:0] comp720minVal;
    wire [5:0] comp720minI, comp720minJ;
    Comparator comp720(SADValues[557*12 +: 12], 8, 45, SADValues[620*12 +: 12], 9, 44, comp720minVal, comp720minI, comp720minJ);
    wire [11:0] comp721minVal;
    wire [5:0] comp721minI, comp721minJ;
    Comparator comp721(SADValues[683*12 +: 12], 10, 43, SADValues[746*12 +: 12], 11, 42, comp721minVal, comp721minI, comp721minJ);
    wire [11:0] comp722minVal;
    wire [5:0] comp722minI, comp722minJ;
    Comparator comp722(SADValues[809*12 +: 12], 12, 41, SADValues[872*12 +: 12], 13, 40, comp722minVal, comp722minI, comp722minJ);
    wire [11:0] comp723minVal;
    wire [5:0] comp723minI, comp723minJ;
    Comparator comp723(SADValues[935*12 +: 12], 14, 39, SADValues[998*12 +: 12], 15, 38, comp723minVal, comp723minI, comp723minJ);
    wire [11:0] comp724minVal;
    wire [5:0] comp724minI, comp724minJ;
    Comparator comp724(SADValues[1061*12 +: 12], 16, 37, SADValues[1124*12 +: 12], 17, 36, comp724minVal, comp724minI, comp724minJ);
    wire [11:0] comp725minVal;
    wire [5:0] comp725minI, comp725minJ;
    Comparator comp725(SADValues[1187*12 +: 12], 18, 35, SADValues[1250*12 +: 12], 19, 34, comp725minVal, comp725minI, comp725minJ);
    wire [11:0] comp726minVal;
    wire [5:0] comp726minI, comp726minJ;
    Comparator comp726(SADValues[1313*12 +: 12], 20, 33, SADValues[1376*12 +: 12], 21, 32, comp726minVal, comp726minI, comp726minJ);
    wire [11:0] comp727minVal;
    wire [5:0] comp727minI, comp727minJ;
    Comparator comp727(SADValues[1439*12 +: 12], 22, 31, SADValues[1502*12 +: 12], 23, 30, comp727minVal, comp727minI, comp727minJ);
    wire [11:0] comp728minVal;
    wire [5:0] comp728minI, comp728minJ;
    Comparator comp728(SADValues[1565*12 +: 12], 24, 29, SADValues[1628*12 +: 12], 25, 28, comp728minVal, comp728minI, comp728minJ);
    wire [11:0] comp729minVal;
    wire [5:0] comp729minI, comp729minJ;
    Comparator comp729(SADValues[1691*12 +: 12], 26, 27, SADValues[1754*12 +: 12], 27, 26, comp729minVal, comp729minI, comp729minJ);
    wire [11:0] comp730minVal;
    wire [5:0] comp730minI, comp730minJ;
    Comparator comp730(SADValues[1817*12 +: 12], 28, 25, SADValues[1880*12 +: 12], 29, 24, comp730minVal, comp730minI, comp730minJ);
    wire [11:0] comp731minVal;
    wire [5:0] comp731minI, comp731minJ;
    Comparator comp731(SADValues[1943*12 +: 12], 30, 23, SADValues[2006*12 +: 12], 31, 22, comp731minVal, comp731minI, comp731minJ);
    wire [11:0] comp732minVal;
    wire [5:0] comp732minI, comp732minJ;
    Comparator comp732(SADValues[2069*12 +: 12], 32, 21, SADValues[2132*12 +: 12], 33, 20, comp732minVal, comp732minI, comp732minJ);
    wire [11:0] comp733minVal;
    wire [5:0] comp733minI, comp733minJ;
    Comparator comp733(SADValues[2195*12 +: 12], 34, 19, SADValues[2258*12 +: 12], 35, 18, comp733minVal, comp733minI, comp733minJ);
    wire [11:0] comp734minVal;
    wire [5:0] comp734minI, comp734minJ;
    Comparator comp734(SADValues[2321*12 +: 12], 36, 17, SADValues[2384*12 +: 12], 37, 16, comp734minVal, comp734minI, comp734minJ);
    wire [11:0] comp735minVal;
    wire [5:0] comp735minI, comp735minJ;
    Comparator comp735(SADValues[2447*12 +: 12], 38, 15, SADValues[2510*12 +: 12], 39, 14, comp735minVal, comp735minI, comp735minJ);
    wire [11:0] comp736minVal;
    wire [5:0] comp736minI, comp736minJ;
    Comparator comp736(SADValues[2573*12 +: 12], 40, 13, SADValues[2636*12 +: 12], 41, 12, comp736minVal, comp736minI, comp736minJ);
    wire [11:0] comp737minVal;
    wire [5:0] comp737minI, comp737minJ;
    Comparator comp737(SADValues[2699*12 +: 12], 42, 11, SADValues[2762*12 +: 12], 43, 10, comp737minVal, comp737minI, comp737minJ);
    wire [11:0] comp738minVal;
    wire [5:0] comp738minI, comp738minJ;
    Comparator comp738(SADValues[2825*12 +: 12], 44, 9, SADValues[2888*12 +: 12], 45, 8, comp738minVal, comp738minI, comp738minJ);
    wire [11:0] comp739minVal;
    wire [5:0] comp739minI, comp739minJ;
    Comparator comp739(SADValues[2951*12 +: 12], 46, 7, SADValues[3014*12 +: 12], 47, 6, comp739minVal, comp739minI, comp739minJ);
    wire [11:0] comp740minVal;
    wire [5:0] comp740minI, comp740minJ;
    Comparator comp740(SADValues[3077*12 +: 12], 48, 5, SADValues[3140*12 +: 12], 49, 4, comp740minVal, comp740minI, comp740minJ);
    wire [11:0] comp741minVal;
    wire [5:0] comp741minI, comp741minJ;
    Comparator comp741(SADValues[3203*12 +: 12], 50, 3, SADValues[3266*12 +: 12], 51, 2, comp741minVal, comp741minI, comp741minJ);
    wire [11:0] comp742minVal;
    wire [5:0] comp742minI, comp742minJ;
    Comparator comp742(SADValues[3329*12 +: 12], 52, 1, SADValues[3392*12 +: 12], 53, 0, comp742minVal, comp742minI, comp742minJ);
    wire [11:0] comp743minVal;
    wire [5:0] comp743minI, comp743minJ;
    Comparator comp743(SADValues[3456*12 +: 12], 54, 0, SADValues[3393*12 +: 12], 53, 1, comp743minVal, comp743minI, comp743minJ);
    wire [11:0] comp744minVal;
    wire [5:0] comp744minI, comp744minJ;
    Comparator comp744(SADValues[3330*12 +: 12], 52, 2, SADValues[3267*12 +: 12], 51, 3, comp744minVal, comp744minI, comp744minJ);
    wire [11:0] comp745minVal;
    wire [5:0] comp745minI, comp745minJ;
    Comparator comp745(SADValues[3204*12 +: 12], 50, 4, SADValues[3141*12 +: 12], 49, 5, comp745minVal, comp745minI, comp745minJ);
    wire [11:0] comp746minVal;
    wire [5:0] comp746minI, comp746minJ;
    Comparator comp746(SADValues[3078*12 +: 12], 48, 6, SADValues[3015*12 +: 12], 47, 7, comp746minVal, comp746minI, comp746minJ);
    wire [11:0] comp747minVal;
    wire [5:0] comp747minI, comp747minJ;
    Comparator comp747(SADValues[2952*12 +: 12], 46, 8, SADValues[2889*12 +: 12], 45, 9, comp747minVal, comp747minI, comp747minJ);
    wire [11:0] comp748minVal;
    wire [5:0] comp748minI, comp748minJ;
    Comparator comp748(SADValues[2826*12 +: 12], 44, 10, SADValues[2763*12 +: 12], 43, 11, comp748minVal, comp748minI, comp748minJ);
    wire [11:0] comp749minVal;
    wire [5:0] comp749minI, comp749minJ;
    Comparator comp749(SADValues[2700*12 +: 12], 42, 12, SADValues[2637*12 +: 12], 41, 13, comp749minVal, comp749minI, comp749minJ);
    wire [11:0] comp750minVal;
    wire [5:0] comp750minI, comp750minJ;
    Comparator comp750(SADValues[2574*12 +: 12], 40, 14, SADValues[2511*12 +: 12], 39, 15, comp750minVal, comp750minI, comp750minJ);
    wire [11:0] comp751minVal;
    wire [5:0] comp751minI, comp751minJ;
    Comparator comp751(SADValues[2448*12 +: 12], 38, 16, SADValues[2385*12 +: 12], 37, 17, comp751minVal, comp751minI, comp751minJ);
    wire [11:0] comp752minVal;
    wire [5:0] comp752minI, comp752minJ;
    Comparator comp752(SADValues[2322*12 +: 12], 36, 18, SADValues[2259*12 +: 12], 35, 19, comp752minVal, comp752minI, comp752minJ);
    wire [11:0] comp753minVal;
    wire [5:0] comp753minI, comp753minJ;
    Comparator comp753(SADValues[2196*12 +: 12], 34, 20, SADValues[2133*12 +: 12], 33, 21, comp753minVal, comp753minI, comp753minJ);
    wire [11:0] comp754minVal;
    wire [5:0] comp754minI, comp754minJ;
    Comparator comp754(SADValues[2070*12 +: 12], 32, 22, SADValues[2007*12 +: 12], 31, 23, comp754minVal, comp754minI, comp754minJ);
    wire [11:0] comp755minVal;
    wire [5:0] comp755minI, comp755minJ;
    Comparator comp755(SADValues[1944*12 +: 12], 30, 24, SADValues[1881*12 +: 12], 29, 25, comp755minVal, comp755minI, comp755minJ);
    wire [11:0] comp756minVal;
    wire [5:0] comp756minI, comp756minJ;
    Comparator comp756(SADValues[1818*12 +: 12], 28, 26, SADValues[1755*12 +: 12], 27, 27, comp756minVal, comp756minI, comp756minJ);
    wire [11:0] comp757minVal;
    wire [5:0] comp757minI, comp757minJ;
    Comparator comp757(SADValues[1692*12 +: 12], 26, 28, SADValues[1629*12 +: 12], 25, 29, comp757minVal, comp757minI, comp757minJ);
    wire [11:0] comp758minVal;
    wire [5:0] comp758minI, comp758minJ;
    Comparator comp758(SADValues[1566*12 +: 12], 24, 30, SADValues[1503*12 +: 12], 23, 31, comp758minVal, comp758minI, comp758minJ);
    wire [11:0] comp759minVal;
    wire [5:0] comp759minI, comp759minJ;
    Comparator comp759(SADValues[1440*12 +: 12], 22, 32, SADValues[1377*12 +: 12], 21, 33, comp759minVal, comp759minI, comp759minJ);
    wire [11:0] comp760minVal;
    wire [5:0] comp760minI, comp760minJ;
    Comparator comp760(SADValues[1314*12 +: 12], 20, 34, SADValues[1251*12 +: 12], 19, 35, comp760minVal, comp760minI, comp760minJ);
    wire [11:0] comp761minVal;
    wire [5:0] comp761minI, comp761minJ;
    Comparator comp761(SADValues[1188*12 +: 12], 18, 36, SADValues[1125*12 +: 12], 17, 37, comp761minVal, comp761minI, comp761minJ);
    wire [11:0] comp762minVal;
    wire [5:0] comp762minI, comp762minJ;
    Comparator comp762(SADValues[1062*12 +: 12], 16, 38, SADValues[999*12 +: 12], 15, 39, comp762minVal, comp762minI, comp762minJ);
    wire [11:0] comp763minVal;
    wire [5:0] comp763minI, comp763minJ;
    Comparator comp763(SADValues[936*12 +: 12], 14, 40, SADValues[873*12 +: 12], 13, 41, comp763minVal, comp763minI, comp763minJ);
    wire [11:0] comp764minVal;
    wire [5:0] comp764minI, comp764minJ;
    Comparator comp764(SADValues[810*12 +: 12], 12, 42, SADValues[747*12 +: 12], 11, 43, comp764minVal, comp764minI, comp764minJ);
    wire [11:0] comp765minVal;
    wire [5:0] comp765minI, comp765minJ;
    Comparator comp765(SADValues[684*12 +: 12], 10, 44, SADValues[621*12 +: 12], 9, 45, comp765minVal, comp765minI, comp765minJ);
    wire [11:0] comp766minVal;
    wire [5:0] comp766minI, comp766minJ;
    Comparator comp766(SADValues[558*12 +: 12], 8, 46, SADValues[495*12 +: 12], 7, 47, comp766minVal, comp766minI, comp766minJ);
    wire [11:0] comp767minVal;
    wire [5:0] comp767minI, comp767minJ;
    Comparator comp767(SADValues[432*12 +: 12], 6, 48, SADValues[369*12 +: 12], 5, 49, comp767minVal, comp767minI, comp767minJ);
    wire [11:0] comp768minVal;
    wire [5:0] comp768minI, comp768minJ;
    Comparator comp768(SADValues[306*12 +: 12], 4, 50, SADValues[243*12 +: 12], 3, 51, comp768minVal, comp768minI, comp768minJ);
    wire [11:0] comp769minVal;
    wire [5:0] comp769minI, comp769minJ;
    Comparator comp769(SADValues[180*12 +: 12], 2, 52, SADValues[117*12 +: 12], 1, 53, comp769minVal, comp769minI, comp769minJ);
    wire [11:0] comp770minVal;
    wire [5:0] comp770minI, comp770minJ;
    Comparator comp770(SADValues[54*12 +: 12], 0, 54, SADValues[55*12 +: 12], 0, 55, comp770minVal, comp770minI, comp770minJ);
    wire [11:0] comp771minVal;
    wire [5:0] comp771minI, comp771minJ;
    Comparator comp771(SADValues[118*12 +: 12], 1, 54, SADValues[181*12 +: 12], 2, 53, comp771minVal, comp771minI, comp771minJ);
    wire [11:0] comp772minVal;
    wire [5:0] comp772minI, comp772minJ;
    Comparator comp772(SADValues[244*12 +: 12], 3, 52, SADValues[307*12 +: 12], 4, 51, comp772minVal, comp772minI, comp772minJ);
    wire [11:0] comp773minVal;
    wire [5:0] comp773minI, comp773minJ;
    Comparator comp773(SADValues[370*12 +: 12], 5, 50, SADValues[433*12 +: 12], 6, 49, comp773minVal, comp773minI, comp773minJ);
    wire [11:0] comp774minVal;
    wire [5:0] comp774minI, comp774minJ;
    Comparator comp774(SADValues[496*12 +: 12], 7, 48, SADValues[559*12 +: 12], 8, 47, comp774minVal, comp774minI, comp774minJ);
    wire [11:0] comp775minVal;
    wire [5:0] comp775minI, comp775minJ;
    Comparator comp775(SADValues[622*12 +: 12], 9, 46, SADValues[685*12 +: 12], 10, 45, comp775minVal, comp775minI, comp775minJ);
    wire [11:0] comp776minVal;
    wire [5:0] comp776minI, comp776minJ;
    Comparator comp776(SADValues[748*12 +: 12], 11, 44, SADValues[811*12 +: 12], 12, 43, comp776minVal, comp776minI, comp776minJ);
    wire [11:0] comp777minVal;
    wire [5:0] comp777minI, comp777minJ;
    Comparator comp777(SADValues[874*12 +: 12], 13, 42, SADValues[937*12 +: 12], 14, 41, comp777minVal, comp777minI, comp777minJ);
    wire [11:0] comp778minVal;
    wire [5:0] comp778minI, comp778minJ;
    Comparator comp778(SADValues[1000*12 +: 12], 15, 40, SADValues[1063*12 +: 12], 16, 39, comp778minVal, comp778minI, comp778minJ);
    wire [11:0] comp779minVal;
    wire [5:0] comp779minI, comp779minJ;
    Comparator comp779(SADValues[1126*12 +: 12], 17, 38, SADValues[1189*12 +: 12], 18, 37, comp779minVal, comp779minI, comp779minJ);
    wire [11:0] comp780minVal;
    wire [5:0] comp780minI, comp780minJ;
    Comparator comp780(SADValues[1252*12 +: 12], 19, 36, SADValues[1315*12 +: 12], 20, 35, comp780minVal, comp780minI, comp780minJ);
    wire [11:0] comp781minVal;
    wire [5:0] comp781minI, comp781minJ;
    Comparator comp781(SADValues[1378*12 +: 12], 21, 34, SADValues[1441*12 +: 12], 22, 33, comp781minVal, comp781minI, comp781minJ);
    wire [11:0] comp782minVal;
    wire [5:0] comp782minI, comp782minJ;
    Comparator comp782(SADValues[1504*12 +: 12], 23, 32, SADValues[1567*12 +: 12], 24, 31, comp782minVal, comp782minI, comp782minJ);
    wire [11:0] comp783minVal;
    wire [5:0] comp783minI, comp783minJ;
    Comparator comp783(SADValues[1630*12 +: 12], 25, 30, SADValues[1693*12 +: 12], 26, 29, comp783minVal, comp783minI, comp783minJ);
    wire [11:0] comp784minVal;
    wire [5:0] comp784minI, comp784minJ;
    Comparator comp784(SADValues[1756*12 +: 12], 27, 28, SADValues[1819*12 +: 12], 28, 27, comp784minVal, comp784minI, comp784minJ);
    wire [11:0] comp785minVal;
    wire [5:0] comp785minI, comp785minJ;
    Comparator comp785(SADValues[1882*12 +: 12], 29, 26, SADValues[1945*12 +: 12], 30, 25, comp785minVal, comp785minI, comp785minJ);
    wire [11:0] comp786minVal;
    wire [5:0] comp786minI, comp786minJ;
    Comparator comp786(SADValues[2008*12 +: 12], 31, 24, SADValues[2071*12 +: 12], 32, 23, comp786minVal, comp786minI, comp786minJ);
    wire [11:0] comp787minVal;
    wire [5:0] comp787minI, comp787minJ;
    Comparator comp787(SADValues[2134*12 +: 12], 33, 22, SADValues[2197*12 +: 12], 34, 21, comp787minVal, comp787minI, comp787minJ);
    wire [11:0] comp788minVal;
    wire [5:0] comp788minI, comp788minJ;
    Comparator comp788(SADValues[2260*12 +: 12], 35, 20, SADValues[2323*12 +: 12], 36, 19, comp788minVal, comp788minI, comp788minJ);
    wire [11:0] comp789minVal;
    wire [5:0] comp789minI, comp789minJ;
    Comparator comp789(SADValues[2386*12 +: 12], 37, 18, SADValues[2449*12 +: 12], 38, 17, comp789minVal, comp789minI, comp789minJ);
    wire [11:0] comp790minVal;
    wire [5:0] comp790minI, comp790minJ;
    Comparator comp790(SADValues[2512*12 +: 12], 39, 16, SADValues[2575*12 +: 12], 40, 15, comp790minVal, comp790minI, comp790minJ);
    wire [11:0] comp791minVal;
    wire [5:0] comp791minI, comp791minJ;
    Comparator comp791(SADValues[2638*12 +: 12], 41, 14, SADValues[2701*12 +: 12], 42, 13, comp791minVal, comp791minI, comp791minJ);
    wire [11:0] comp792minVal;
    wire [5:0] comp792minI, comp792minJ;
    Comparator comp792(SADValues[2764*12 +: 12], 43, 12, SADValues[2827*12 +: 12], 44, 11, comp792minVal, comp792minI, comp792minJ);
    wire [11:0] comp793minVal;
    wire [5:0] comp793minI, comp793minJ;
    Comparator comp793(SADValues[2890*12 +: 12], 45, 10, SADValues[2953*12 +: 12], 46, 9, comp793minVal, comp793minI, comp793minJ);
    wire [11:0] comp794minVal;
    wire [5:0] comp794minI, comp794minJ;
    Comparator comp794(SADValues[3016*12 +: 12], 47, 8, SADValues[3079*12 +: 12], 48, 7, comp794minVal, comp794minI, comp794minJ);
    wire [11:0] comp795minVal;
    wire [5:0] comp795minI, comp795minJ;
    Comparator comp795(SADValues[3142*12 +: 12], 49, 6, SADValues[3205*12 +: 12], 50, 5, comp795minVal, comp795minI, comp795minJ);
    wire [11:0] comp796minVal;
    wire [5:0] comp796minI, comp796minJ;
    Comparator comp796(SADValues[3268*12 +: 12], 51, 4, SADValues[3331*12 +: 12], 52, 3, comp796minVal, comp796minI, comp796minJ);
    wire [11:0] comp797minVal;
    wire [5:0] comp797minI, comp797minJ;
    Comparator comp797(SADValues[3394*12 +: 12], 53, 2, SADValues[3457*12 +: 12], 54, 1, comp797minVal, comp797minI, comp797minJ);
    wire [11:0] comp798minVal;
    wire [5:0] comp798minI, comp798minJ;
    Comparator comp798(SADValues[3520*12 +: 12], 55, 0, SADValues[3584*12 +: 12], 56, 0, comp798minVal, comp798minI, comp798minJ);
    wire [11:0] comp799minVal;
    wire [5:0] comp799minI, comp799minJ;
    Comparator comp799(SADValues[3521*12 +: 12], 55, 1, SADValues[3458*12 +: 12], 54, 2, comp799minVal, comp799minI, comp799minJ);
    wire [11:0] comp800minVal;
    wire [5:0] comp800minI, comp800minJ;
    Comparator comp800(SADValues[3395*12 +: 12], 53, 3, SADValues[3332*12 +: 12], 52, 4, comp800minVal, comp800minI, comp800minJ);
    wire [11:0] comp801minVal;
    wire [5:0] comp801minI, comp801minJ;
    Comparator comp801(SADValues[3269*12 +: 12], 51, 5, SADValues[3206*12 +: 12], 50, 6, comp801minVal, comp801minI, comp801minJ);
    wire [11:0] comp802minVal;
    wire [5:0] comp802minI, comp802minJ;
    Comparator comp802(SADValues[3143*12 +: 12], 49, 7, SADValues[3080*12 +: 12], 48, 8, comp802minVal, comp802minI, comp802minJ);
    wire [11:0] comp803minVal;
    wire [5:0] comp803minI, comp803minJ;
    Comparator comp803(SADValues[3017*12 +: 12], 47, 9, SADValues[2954*12 +: 12], 46, 10, comp803minVal, comp803minI, comp803minJ);
    wire [11:0] comp804minVal;
    wire [5:0] comp804minI, comp804minJ;
    Comparator comp804(SADValues[2891*12 +: 12], 45, 11, SADValues[2828*12 +: 12], 44, 12, comp804minVal, comp804minI, comp804minJ);
    wire [11:0] comp805minVal;
    wire [5:0] comp805minI, comp805minJ;
    Comparator comp805(SADValues[2765*12 +: 12], 43, 13, SADValues[2702*12 +: 12], 42, 14, comp805minVal, comp805minI, comp805minJ);
    wire [11:0] comp806minVal;
    wire [5:0] comp806minI, comp806minJ;
    Comparator comp806(SADValues[2639*12 +: 12], 41, 15, SADValues[2576*12 +: 12], 40, 16, comp806minVal, comp806minI, comp806minJ);
    wire [11:0] comp807minVal;
    wire [5:0] comp807minI, comp807minJ;
    Comparator comp807(SADValues[2513*12 +: 12], 39, 17, SADValues[2450*12 +: 12], 38, 18, comp807minVal, comp807minI, comp807minJ);
    wire [11:0] comp808minVal;
    wire [5:0] comp808minI, comp808minJ;
    Comparator comp808(SADValues[2387*12 +: 12], 37, 19, SADValues[2324*12 +: 12], 36, 20, comp808minVal, comp808minI, comp808minJ);
    wire [11:0] comp809minVal;
    wire [5:0] comp809minI, comp809minJ;
    Comparator comp809(SADValues[2261*12 +: 12], 35, 21, SADValues[2198*12 +: 12], 34, 22, comp809minVal, comp809minI, comp809minJ);
    wire [11:0] comp810minVal;
    wire [5:0] comp810minI, comp810minJ;
    Comparator comp810(SADValues[2135*12 +: 12], 33, 23, SADValues[2072*12 +: 12], 32, 24, comp810minVal, comp810minI, comp810minJ);
    wire [11:0] comp811minVal;
    wire [5:0] comp811minI, comp811minJ;
    Comparator comp811(SADValues[2009*12 +: 12], 31, 25, SADValues[1946*12 +: 12], 30, 26, comp811minVal, comp811minI, comp811minJ);
    wire [11:0] comp812minVal;
    wire [5:0] comp812minI, comp812minJ;
    Comparator comp812(SADValues[1883*12 +: 12], 29, 27, SADValues[1820*12 +: 12], 28, 28, comp812minVal, comp812minI, comp812minJ);
    wire [11:0] comp813minVal;
    wire [5:0] comp813minI, comp813minJ;
    Comparator comp813(SADValues[1757*12 +: 12], 27, 29, SADValues[1694*12 +: 12], 26, 30, comp813minVal, comp813minI, comp813minJ);
    wire [11:0] comp814minVal;
    wire [5:0] comp814minI, comp814minJ;
    Comparator comp814(SADValues[1631*12 +: 12], 25, 31, SADValues[1568*12 +: 12], 24, 32, comp814minVal, comp814minI, comp814minJ);
    wire [11:0] comp815minVal;
    wire [5:0] comp815minI, comp815minJ;
    Comparator comp815(SADValues[1505*12 +: 12], 23, 33, SADValues[1442*12 +: 12], 22, 34, comp815minVal, comp815minI, comp815minJ);
    wire [11:0] comp816minVal;
    wire [5:0] comp816minI, comp816minJ;
    Comparator comp816(SADValues[1379*12 +: 12], 21, 35, SADValues[1316*12 +: 12], 20, 36, comp816minVal, comp816minI, comp816minJ);
    wire [11:0] comp817minVal;
    wire [5:0] comp817minI, comp817minJ;
    Comparator comp817(SADValues[1253*12 +: 12], 19, 37, SADValues[1190*12 +: 12], 18, 38, comp817minVal, comp817minI, comp817minJ);
    wire [11:0] comp818minVal;
    wire [5:0] comp818minI, comp818minJ;
    Comparator comp818(SADValues[1127*12 +: 12], 17, 39, SADValues[1064*12 +: 12], 16, 40, comp818minVal, comp818minI, comp818minJ);
    wire [11:0] comp819minVal;
    wire [5:0] comp819minI, comp819minJ;
    Comparator comp819(SADValues[1001*12 +: 12], 15, 41, SADValues[938*12 +: 12], 14, 42, comp819minVal, comp819minI, comp819minJ);
    wire [11:0] comp820minVal;
    wire [5:0] comp820minI, comp820minJ;
    Comparator comp820(SADValues[875*12 +: 12], 13, 43, SADValues[812*12 +: 12], 12, 44, comp820minVal, comp820minI, comp820minJ);
    wire [11:0] comp821minVal;
    wire [5:0] comp821minI, comp821minJ;
    Comparator comp821(SADValues[749*12 +: 12], 11, 45, SADValues[686*12 +: 12], 10, 46, comp821minVal, comp821minI, comp821minJ);
    wire [11:0] comp822minVal;
    wire [5:0] comp822minI, comp822minJ;
    Comparator comp822(SADValues[623*12 +: 12], 9, 47, SADValues[560*12 +: 12], 8, 48, comp822minVal, comp822minI, comp822minJ);
    wire [11:0] comp823minVal;
    wire [5:0] comp823minI, comp823minJ;
    Comparator comp823(SADValues[497*12 +: 12], 7, 49, SADValues[434*12 +: 12], 6, 50, comp823minVal, comp823minI, comp823minJ);
    wire [11:0] comp824minVal;
    wire [5:0] comp824minI, comp824minJ;
    Comparator comp824(SADValues[371*12 +: 12], 5, 51, SADValues[308*12 +: 12], 4, 52, comp824minVal, comp824minI, comp824minJ);
    wire [11:0] comp825minVal;
    wire [5:0] comp825minI, comp825minJ;
    Comparator comp825(SADValues[245*12 +: 12], 3, 53, SADValues[182*12 +: 12], 2, 54, comp825minVal, comp825minI, comp825minJ);
    wire [11:0] comp826minVal;
    wire [5:0] comp826minI, comp826minJ;
    Comparator comp826(SADValues[119*12 +: 12], 1, 55, SADValues[56*12 +: 12], 0, 56, comp826minVal, comp826minI, comp826minJ);
    wire [11:0] comp827minVal;
    wire [5:0] comp827minI, comp827minJ;
    Comparator comp827(SADValues[57*12 +: 12], 0, 57, SADValues[120*12 +: 12], 1, 56, comp827minVal, comp827minI, comp827minJ);
    wire [11:0] comp828minVal;
    wire [5:0] comp828minI, comp828minJ;
    Comparator comp828(SADValues[183*12 +: 12], 2, 55, SADValues[246*12 +: 12], 3, 54, comp828minVal, comp828minI, comp828minJ);
    wire [11:0] comp829minVal;
    wire [5:0] comp829minI, comp829minJ;
    Comparator comp829(SADValues[309*12 +: 12], 4, 53, SADValues[372*12 +: 12], 5, 52, comp829minVal, comp829minI, comp829minJ);
    wire [11:0] comp830minVal;
    wire [5:0] comp830minI, comp830minJ;
    Comparator comp830(SADValues[435*12 +: 12], 6, 51, SADValues[498*12 +: 12], 7, 50, comp830minVal, comp830minI, comp830minJ);
    wire [11:0] comp831minVal;
    wire [5:0] comp831minI, comp831minJ;
    Comparator comp831(SADValues[561*12 +: 12], 8, 49, SADValues[624*12 +: 12], 9, 48, comp831minVal, comp831minI, comp831minJ);
    wire [11:0] comp832minVal;
    wire [5:0] comp832minI, comp832minJ;
    Comparator comp832(SADValues[687*12 +: 12], 10, 47, SADValues[750*12 +: 12], 11, 46, comp832minVal, comp832minI, comp832minJ);
    wire [11:0] comp833minVal;
    wire [5:0] comp833minI, comp833minJ;
    Comparator comp833(SADValues[813*12 +: 12], 12, 45, SADValues[876*12 +: 12], 13, 44, comp833minVal, comp833minI, comp833minJ);
    wire [11:0] comp834minVal;
    wire [5:0] comp834minI, comp834minJ;
    Comparator comp834(SADValues[939*12 +: 12], 14, 43, SADValues[1002*12 +: 12], 15, 42, comp834minVal, comp834minI, comp834minJ);
    wire [11:0] comp835minVal;
    wire [5:0] comp835minI, comp835minJ;
    Comparator comp835(SADValues[1065*12 +: 12], 16, 41, SADValues[1128*12 +: 12], 17, 40, comp835minVal, comp835minI, comp835minJ);
    wire [11:0] comp836minVal;
    wire [5:0] comp836minI, comp836minJ;
    Comparator comp836(SADValues[1191*12 +: 12], 18, 39, SADValues[1254*12 +: 12], 19, 38, comp836minVal, comp836minI, comp836minJ);
    wire [11:0] comp837minVal;
    wire [5:0] comp837minI, comp837minJ;
    Comparator comp837(SADValues[1317*12 +: 12], 20, 37, SADValues[1380*12 +: 12], 21, 36, comp837minVal, comp837minI, comp837minJ);
    wire [11:0] comp838minVal;
    wire [5:0] comp838minI, comp838minJ;
    Comparator comp838(SADValues[1443*12 +: 12], 22, 35, SADValues[1506*12 +: 12], 23, 34, comp838minVal, comp838minI, comp838minJ);
    wire [11:0] comp839minVal;
    wire [5:0] comp839minI, comp839minJ;
    Comparator comp839(SADValues[1569*12 +: 12], 24, 33, SADValues[1632*12 +: 12], 25, 32, comp839minVal, comp839minI, comp839minJ);
    wire [11:0] comp840minVal;
    wire [5:0] comp840minI, comp840minJ;
    Comparator comp840(SADValues[1695*12 +: 12], 26, 31, SADValues[1758*12 +: 12], 27, 30, comp840minVal, comp840minI, comp840minJ);
    wire [11:0] comp841minVal;
    wire [5:0] comp841minI, comp841minJ;
    Comparator comp841(SADValues[1821*12 +: 12], 28, 29, SADValues[1884*12 +: 12], 29, 28, comp841minVal, comp841minI, comp841minJ);
    wire [11:0] comp842minVal;
    wire [5:0] comp842minI, comp842minJ;
    Comparator comp842(SADValues[1947*12 +: 12], 30, 27, SADValues[2010*12 +: 12], 31, 26, comp842minVal, comp842minI, comp842minJ);
    wire [11:0] comp843minVal;
    wire [5:0] comp843minI, comp843minJ;
    Comparator comp843(SADValues[2073*12 +: 12], 32, 25, SADValues[2136*12 +: 12], 33, 24, comp843minVal, comp843minI, comp843minJ);
    wire [11:0] comp844minVal;
    wire [5:0] comp844minI, comp844minJ;
    Comparator comp844(SADValues[2199*12 +: 12], 34, 23, SADValues[2262*12 +: 12], 35, 22, comp844minVal, comp844minI, comp844minJ);
    wire [11:0] comp845minVal;
    wire [5:0] comp845minI, comp845minJ;
    Comparator comp845(SADValues[2325*12 +: 12], 36, 21, SADValues[2388*12 +: 12], 37, 20, comp845minVal, comp845minI, comp845minJ);
    wire [11:0] comp846minVal;
    wire [5:0] comp846minI, comp846minJ;
    Comparator comp846(SADValues[2451*12 +: 12], 38, 19, SADValues[2514*12 +: 12], 39, 18, comp846minVal, comp846minI, comp846minJ);
    wire [11:0] comp847minVal;
    wire [5:0] comp847minI, comp847minJ;
    Comparator comp847(SADValues[2577*12 +: 12], 40, 17, SADValues[2640*12 +: 12], 41, 16, comp847minVal, comp847minI, comp847minJ);
    wire [11:0] comp848minVal;
    wire [5:0] comp848minI, comp848minJ;
    Comparator comp848(SADValues[2703*12 +: 12], 42, 15, SADValues[2766*12 +: 12], 43, 14, comp848minVal, comp848minI, comp848minJ);
    wire [11:0] comp849minVal;
    wire [5:0] comp849minI, comp849minJ;
    Comparator comp849(SADValues[2829*12 +: 12], 44, 13, SADValues[2892*12 +: 12], 45, 12, comp849minVal, comp849minI, comp849minJ);
    wire [11:0] comp850minVal;
    wire [5:0] comp850minI, comp850minJ;
    Comparator comp850(SADValues[2955*12 +: 12], 46, 11, SADValues[3018*12 +: 12], 47, 10, comp850minVal, comp850minI, comp850minJ);
    wire [11:0] comp851minVal;
    wire [5:0] comp851minI, comp851minJ;
    Comparator comp851(SADValues[3081*12 +: 12], 48, 9, SADValues[3144*12 +: 12], 49, 8, comp851minVal, comp851minI, comp851minJ);
    wire [11:0] comp852minVal;
    wire [5:0] comp852minI, comp852minJ;
    Comparator comp852(SADValues[3207*12 +: 12], 50, 7, SADValues[3270*12 +: 12], 51, 6, comp852minVal, comp852minI, comp852minJ);
    wire [11:0] comp853minVal;
    wire [5:0] comp853minI, comp853minJ;
    Comparator comp853(SADValues[3333*12 +: 12], 52, 5, SADValues[3396*12 +: 12], 53, 4, comp853minVal, comp853minI, comp853minJ);
    wire [11:0] comp854minVal;
    wire [5:0] comp854minI, comp854minJ;
    Comparator comp854(SADValues[3459*12 +: 12], 54, 3, SADValues[3522*12 +: 12], 55, 2, comp854minVal, comp854minI, comp854minJ);
    wire [11:0] comp855minVal;
    wire [5:0] comp855minI, comp855minJ;
    Comparator comp855(SADValues[3585*12 +: 12], 56, 1, SADValues[3648*12 +: 12], 57, 0, comp855minVal, comp855minI, comp855minJ);
    wire [11:0] comp856minVal;
    wire [5:0] comp856minI, comp856minJ;
    Comparator comp856(SADValues[3712*12 +: 12], 58, 0, SADValues[3649*12 +: 12], 57, 1, comp856minVal, comp856minI, comp856minJ);
    wire [11:0] comp857minVal;
    wire [5:0] comp857minI, comp857minJ;
    Comparator comp857(SADValues[3586*12 +: 12], 56, 2, SADValues[3523*12 +: 12], 55, 3, comp857minVal, comp857minI, comp857minJ);
    wire [11:0] comp858minVal;
    wire [5:0] comp858minI, comp858minJ;
    Comparator comp858(SADValues[3460*12 +: 12], 54, 4, SADValues[3397*12 +: 12], 53, 5, comp858minVal, comp858minI, comp858minJ);
    wire [11:0] comp859minVal;
    wire [5:0] comp859minI, comp859minJ;
    Comparator comp859(SADValues[3334*12 +: 12], 52, 6, SADValues[3271*12 +: 12], 51, 7, comp859minVal, comp859minI, comp859minJ);
    wire [11:0] comp860minVal;
    wire [5:0] comp860minI, comp860minJ;
    Comparator comp860(SADValues[3208*12 +: 12], 50, 8, SADValues[3145*12 +: 12], 49, 9, comp860minVal, comp860minI, comp860minJ);
    wire [11:0] comp861minVal;
    wire [5:0] comp861minI, comp861minJ;
    Comparator comp861(SADValues[3082*12 +: 12], 48, 10, SADValues[3019*12 +: 12], 47, 11, comp861minVal, comp861minI, comp861minJ);
    wire [11:0] comp862minVal;
    wire [5:0] comp862minI, comp862minJ;
    Comparator comp862(SADValues[2956*12 +: 12], 46, 12, SADValues[2893*12 +: 12], 45, 13, comp862minVal, comp862minI, comp862minJ);
    wire [11:0] comp863minVal;
    wire [5:0] comp863minI, comp863minJ;
    Comparator comp863(SADValues[2830*12 +: 12], 44, 14, SADValues[2767*12 +: 12], 43, 15, comp863minVal, comp863minI, comp863minJ);
    wire [11:0] comp864minVal;
    wire [5:0] comp864minI, comp864minJ;
    Comparator comp864(SADValues[2704*12 +: 12], 42, 16, SADValues[2641*12 +: 12], 41, 17, comp864minVal, comp864minI, comp864minJ);
    wire [11:0] comp865minVal;
    wire [5:0] comp865minI, comp865minJ;
    Comparator comp865(SADValues[2578*12 +: 12], 40, 18, SADValues[2515*12 +: 12], 39, 19, comp865minVal, comp865minI, comp865minJ);
    wire [11:0] comp866minVal;
    wire [5:0] comp866minI, comp866minJ;
    Comparator comp866(SADValues[2452*12 +: 12], 38, 20, SADValues[2389*12 +: 12], 37, 21, comp866minVal, comp866minI, comp866minJ);
    wire [11:0] comp867minVal;
    wire [5:0] comp867minI, comp867minJ;
    Comparator comp867(SADValues[2326*12 +: 12], 36, 22, SADValues[2263*12 +: 12], 35, 23, comp867minVal, comp867minI, comp867minJ);
    wire [11:0] comp868minVal;
    wire [5:0] comp868minI, comp868minJ;
    Comparator comp868(SADValues[2200*12 +: 12], 34, 24, SADValues[2137*12 +: 12], 33, 25, comp868minVal, comp868minI, comp868minJ);
    wire [11:0] comp869minVal;
    wire [5:0] comp869minI, comp869minJ;
    Comparator comp869(SADValues[2074*12 +: 12], 32, 26, SADValues[2011*12 +: 12], 31, 27, comp869minVal, comp869minI, comp869minJ);
    wire [11:0] comp870minVal;
    wire [5:0] comp870minI, comp870minJ;
    Comparator comp870(SADValues[1948*12 +: 12], 30, 28, SADValues[1885*12 +: 12], 29, 29, comp870minVal, comp870minI, comp870minJ);
    wire [11:0] comp871minVal;
    wire [5:0] comp871minI, comp871minJ;
    Comparator comp871(SADValues[1822*12 +: 12], 28, 30, SADValues[1759*12 +: 12], 27, 31, comp871minVal, comp871minI, comp871minJ);
    wire [11:0] comp872minVal;
    wire [5:0] comp872minI, comp872minJ;
    Comparator comp872(SADValues[1696*12 +: 12], 26, 32, SADValues[1633*12 +: 12], 25, 33, comp872minVal, comp872minI, comp872minJ);
    wire [11:0] comp873minVal;
    wire [5:0] comp873minI, comp873minJ;
    Comparator comp873(SADValues[1570*12 +: 12], 24, 34, SADValues[1507*12 +: 12], 23, 35, comp873minVal, comp873minI, comp873minJ);
    wire [11:0] comp874minVal;
    wire [5:0] comp874minI, comp874minJ;
    Comparator comp874(SADValues[1444*12 +: 12], 22, 36, SADValues[1381*12 +: 12], 21, 37, comp874minVal, comp874minI, comp874minJ);
    wire [11:0] comp875minVal;
    wire [5:0] comp875minI, comp875minJ;
    Comparator comp875(SADValues[1318*12 +: 12], 20, 38, SADValues[1255*12 +: 12], 19, 39, comp875minVal, comp875minI, comp875minJ);
    wire [11:0] comp876minVal;
    wire [5:0] comp876minI, comp876minJ;
    Comparator comp876(SADValues[1192*12 +: 12], 18, 40, SADValues[1129*12 +: 12], 17, 41, comp876minVal, comp876minI, comp876minJ);
    wire [11:0] comp877minVal;
    wire [5:0] comp877minI, comp877minJ;
    Comparator comp877(SADValues[1066*12 +: 12], 16, 42, SADValues[1003*12 +: 12], 15, 43, comp877minVal, comp877minI, comp877minJ);
    wire [11:0] comp878minVal;
    wire [5:0] comp878minI, comp878minJ;
    Comparator comp878(SADValues[940*12 +: 12], 14, 44, SADValues[877*12 +: 12], 13, 45, comp878minVal, comp878minI, comp878minJ);
    wire [11:0] comp879minVal;
    wire [5:0] comp879minI, comp879minJ;
    Comparator comp879(SADValues[814*12 +: 12], 12, 46, SADValues[751*12 +: 12], 11, 47, comp879minVal, comp879minI, comp879minJ);
    wire [11:0] comp880minVal;
    wire [5:0] comp880minI, comp880minJ;
    Comparator comp880(SADValues[688*12 +: 12], 10, 48, SADValues[625*12 +: 12], 9, 49, comp880minVal, comp880minI, comp880minJ);
    wire [11:0] comp881minVal;
    wire [5:0] comp881minI, comp881minJ;
    Comparator comp881(SADValues[562*12 +: 12], 8, 50, SADValues[499*12 +: 12], 7, 51, comp881minVal, comp881minI, comp881minJ);
    wire [11:0] comp882minVal;
    wire [5:0] comp882minI, comp882minJ;
    Comparator comp882(SADValues[436*12 +: 12], 6, 52, SADValues[373*12 +: 12], 5, 53, comp882minVal, comp882minI, comp882minJ);
    wire [11:0] comp883minVal;
    wire [5:0] comp883minI, comp883minJ;
    Comparator comp883(SADValues[310*12 +: 12], 4, 54, SADValues[247*12 +: 12], 3, 55, comp883minVal, comp883minI, comp883minJ);
    wire [11:0] comp884minVal;
    wire [5:0] comp884minI, comp884minJ;
    Comparator comp884(SADValues[184*12 +: 12], 2, 56, SADValues[121*12 +: 12], 1, 57, comp884minVal, comp884minI, comp884minJ);
    wire [11:0] comp885minVal;
    wire [5:0] comp885minI, comp885minJ;
    Comparator comp885(SADValues[58*12 +: 12], 0, 58, SADValues[59*12 +: 12], 0, 59, comp885minVal, comp885minI, comp885minJ);
    wire [11:0] comp886minVal;
    wire [5:0] comp886minI, comp886minJ;
    Comparator comp886(SADValues[122*12 +: 12], 1, 58, SADValues[185*12 +: 12], 2, 57, comp886minVal, comp886minI, comp886minJ);
    wire [11:0] comp887minVal;
    wire [5:0] comp887minI, comp887minJ;
    Comparator comp887(SADValues[248*12 +: 12], 3, 56, SADValues[311*12 +: 12], 4, 55, comp887minVal, comp887minI, comp887minJ);
    wire [11:0] comp888minVal;
    wire [5:0] comp888minI, comp888minJ;
    Comparator comp888(SADValues[374*12 +: 12], 5, 54, SADValues[437*12 +: 12], 6, 53, comp888minVal, comp888minI, comp888minJ);
    wire [11:0] comp889minVal;
    wire [5:0] comp889minI, comp889minJ;
    Comparator comp889(SADValues[500*12 +: 12], 7, 52, SADValues[563*12 +: 12], 8, 51, comp889minVal, comp889minI, comp889minJ);
    wire [11:0] comp890minVal;
    wire [5:0] comp890minI, comp890minJ;
    Comparator comp890(SADValues[626*12 +: 12], 9, 50, SADValues[689*12 +: 12], 10, 49, comp890minVal, comp890minI, comp890minJ);
    wire [11:0] comp891minVal;
    wire [5:0] comp891minI, comp891minJ;
    Comparator comp891(SADValues[752*12 +: 12], 11, 48, SADValues[815*12 +: 12], 12, 47, comp891minVal, comp891minI, comp891minJ);
    wire [11:0] comp892minVal;
    wire [5:0] comp892minI, comp892minJ;
    Comparator comp892(SADValues[878*12 +: 12], 13, 46, SADValues[941*12 +: 12], 14, 45, comp892minVal, comp892minI, comp892minJ);
    wire [11:0] comp893minVal;
    wire [5:0] comp893minI, comp893minJ;
    Comparator comp893(SADValues[1004*12 +: 12], 15, 44, SADValues[1067*12 +: 12], 16, 43, comp893minVal, comp893minI, comp893minJ);
    wire [11:0] comp894minVal;
    wire [5:0] comp894minI, comp894minJ;
    Comparator comp894(SADValues[1130*12 +: 12], 17, 42, SADValues[1193*12 +: 12], 18, 41, comp894minVal, comp894minI, comp894minJ);
    wire [11:0] comp895minVal;
    wire [5:0] comp895minI, comp895minJ;
    Comparator comp895(SADValues[1256*12 +: 12], 19, 40, SADValues[1319*12 +: 12], 20, 39, comp895minVal, comp895minI, comp895minJ);
    wire [11:0] comp896minVal;
    wire [5:0] comp896minI, comp896minJ;
    Comparator comp896(SADValues[1382*12 +: 12], 21, 38, SADValues[1445*12 +: 12], 22, 37, comp896minVal, comp896minI, comp896minJ);
    wire [11:0] comp897minVal;
    wire [5:0] comp897minI, comp897minJ;
    Comparator comp897(SADValues[1508*12 +: 12], 23, 36, SADValues[1571*12 +: 12], 24, 35, comp897minVal, comp897minI, comp897minJ);
    wire [11:0] comp898minVal;
    wire [5:0] comp898minI, comp898minJ;
    Comparator comp898(SADValues[1634*12 +: 12], 25, 34, SADValues[1697*12 +: 12], 26, 33, comp898minVal, comp898minI, comp898minJ);
    wire [11:0] comp899minVal;
    wire [5:0] comp899minI, comp899minJ;
    Comparator comp899(SADValues[1760*12 +: 12], 27, 32, SADValues[1823*12 +: 12], 28, 31, comp899minVal, comp899minI, comp899minJ);
    wire [11:0] comp900minVal;
    wire [5:0] comp900minI, comp900minJ;
    Comparator comp900(SADValues[1886*12 +: 12], 29, 30, SADValues[1949*12 +: 12], 30, 29, comp900minVal, comp900minI, comp900minJ);
    wire [11:0] comp901minVal;
    wire [5:0] comp901minI, comp901minJ;
    Comparator comp901(SADValues[2012*12 +: 12], 31, 28, SADValues[2075*12 +: 12], 32, 27, comp901minVal, comp901minI, comp901minJ);
    wire [11:0] comp902minVal;
    wire [5:0] comp902minI, comp902minJ;
    Comparator comp902(SADValues[2138*12 +: 12], 33, 26, SADValues[2201*12 +: 12], 34, 25, comp902minVal, comp902minI, comp902minJ);
    wire [11:0] comp903minVal;
    wire [5:0] comp903minI, comp903minJ;
    Comparator comp903(SADValues[2264*12 +: 12], 35, 24, SADValues[2327*12 +: 12], 36, 23, comp903minVal, comp903minI, comp903minJ);
    wire [11:0] comp904minVal;
    wire [5:0] comp904minI, comp904minJ;
    Comparator comp904(SADValues[2390*12 +: 12], 37, 22, SADValues[2453*12 +: 12], 38, 21, comp904minVal, comp904minI, comp904minJ);
    wire [11:0] comp905minVal;
    wire [5:0] comp905minI, comp905minJ;
    Comparator comp905(SADValues[2516*12 +: 12], 39, 20, SADValues[2579*12 +: 12], 40, 19, comp905minVal, comp905minI, comp905minJ);
    wire [11:0] comp906minVal;
    wire [5:0] comp906minI, comp906minJ;
    Comparator comp906(SADValues[2642*12 +: 12], 41, 18, SADValues[2705*12 +: 12], 42, 17, comp906minVal, comp906minI, comp906minJ);
    wire [11:0] comp907minVal;
    wire [5:0] comp907minI, comp907minJ;
    Comparator comp907(SADValues[2768*12 +: 12], 43, 16, SADValues[2831*12 +: 12], 44, 15, comp907minVal, comp907minI, comp907minJ);
    wire [11:0] comp908minVal;
    wire [5:0] comp908minI, comp908minJ;
    Comparator comp908(SADValues[2894*12 +: 12], 45, 14, SADValues[2957*12 +: 12], 46, 13, comp908minVal, comp908minI, comp908minJ);
    wire [11:0] comp909minVal;
    wire [5:0] comp909minI, comp909minJ;
    Comparator comp909(SADValues[3020*12 +: 12], 47, 12, SADValues[3083*12 +: 12], 48, 11, comp909minVal, comp909minI, comp909minJ);
    wire [11:0] comp910minVal;
    wire [5:0] comp910minI, comp910minJ;
    Comparator comp910(SADValues[3146*12 +: 12], 49, 10, SADValues[3209*12 +: 12], 50, 9, comp910minVal, comp910minI, comp910minJ);
    wire [11:0] comp911minVal;
    wire [5:0] comp911minI, comp911minJ;
    Comparator comp911(SADValues[3272*12 +: 12], 51, 8, SADValues[3335*12 +: 12], 52, 7, comp911minVal, comp911minI, comp911minJ);
    wire [11:0] comp912minVal;
    wire [5:0] comp912minI, comp912minJ;
    Comparator comp912(SADValues[3398*12 +: 12], 53, 6, SADValues[3461*12 +: 12], 54, 5, comp912minVal, comp912minI, comp912minJ);
    wire [11:0] comp913minVal;
    wire [5:0] comp913minI, comp913minJ;
    Comparator comp913(SADValues[3524*12 +: 12], 55, 4, SADValues[3587*12 +: 12], 56, 3, comp913minVal, comp913minI, comp913minJ);
    wire [11:0] comp914minVal;
    wire [5:0] comp914minI, comp914minJ;
    Comparator comp914(SADValues[3650*12 +: 12], 57, 2, SADValues[3713*12 +: 12], 58, 1, comp914minVal, comp914minI, comp914minJ);
    wire [11:0] comp915minVal;
    wire [5:0] comp915minI, comp915minJ;
    Comparator comp915(SADValues[3776*12 +: 12], 59, 0, SADValues[3840*12 +: 12], 60, 0, comp915minVal, comp915minI, comp915minJ);
    wire [11:0] comp916minVal;
    wire [5:0] comp916minI, comp916minJ;
    Comparator comp916(SADValues[3777*12 +: 12], 59, 1, SADValues[3714*12 +: 12], 58, 2, comp916minVal, comp916minI, comp916minJ);
    wire [11:0] comp917minVal;
    wire [5:0] comp917minI, comp917minJ;
    Comparator comp917(SADValues[3651*12 +: 12], 57, 3, SADValues[3588*12 +: 12], 56, 4, comp917minVal, comp917minI, comp917minJ);
    wire [11:0] comp918minVal;
    wire [5:0] comp918minI, comp918minJ;
    Comparator comp918(SADValues[3525*12 +: 12], 55, 5, SADValues[3462*12 +: 12], 54, 6, comp918minVal, comp918minI, comp918minJ);
    wire [11:0] comp919minVal;
    wire [5:0] comp919minI, comp919minJ;
    Comparator comp919(SADValues[3399*12 +: 12], 53, 7, SADValues[3336*12 +: 12], 52, 8, comp919minVal, comp919minI, comp919minJ);
    wire [11:0] comp920minVal;
    wire [5:0] comp920minI, comp920minJ;
    Comparator comp920(SADValues[3273*12 +: 12], 51, 9, SADValues[3210*12 +: 12], 50, 10, comp920minVal, comp920minI, comp920minJ);
    wire [11:0] comp921minVal;
    wire [5:0] comp921minI, comp921minJ;
    Comparator comp921(SADValues[3147*12 +: 12], 49, 11, SADValues[3084*12 +: 12], 48, 12, comp921minVal, comp921minI, comp921minJ);
    wire [11:0] comp922minVal;
    wire [5:0] comp922minI, comp922minJ;
    Comparator comp922(SADValues[3021*12 +: 12], 47, 13, SADValues[2958*12 +: 12], 46, 14, comp922minVal, comp922minI, comp922minJ);
    wire [11:0] comp923minVal;
    wire [5:0] comp923minI, comp923minJ;
    Comparator comp923(SADValues[2895*12 +: 12], 45, 15, SADValues[2832*12 +: 12], 44, 16, comp923minVal, comp923minI, comp923minJ);
    wire [11:0] comp924minVal;
    wire [5:0] comp924minI, comp924minJ;
    Comparator comp924(SADValues[2769*12 +: 12], 43, 17, SADValues[2706*12 +: 12], 42, 18, comp924minVal, comp924minI, comp924minJ);
    wire [11:0] comp925minVal;
    wire [5:0] comp925minI, comp925minJ;
    Comparator comp925(SADValues[2643*12 +: 12], 41, 19, SADValues[2580*12 +: 12], 40, 20, comp925minVal, comp925minI, comp925minJ);
    wire [11:0] comp926minVal;
    wire [5:0] comp926minI, comp926minJ;
    Comparator comp926(SADValues[2517*12 +: 12], 39, 21, SADValues[2454*12 +: 12], 38, 22, comp926minVal, comp926minI, comp926minJ);
    wire [11:0] comp927minVal;
    wire [5:0] comp927minI, comp927minJ;
    Comparator comp927(SADValues[2391*12 +: 12], 37, 23, SADValues[2328*12 +: 12], 36, 24, comp927minVal, comp927minI, comp927minJ);
    wire [11:0] comp928minVal;
    wire [5:0] comp928minI, comp928minJ;
    Comparator comp928(SADValues[2265*12 +: 12], 35, 25, SADValues[2202*12 +: 12], 34, 26, comp928minVal, comp928minI, comp928minJ);
    wire [11:0] comp929minVal;
    wire [5:0] comp929minI, comp929minJ;
    Comparator comp929(SADValues[2139*12 +: 12], 33, 27, SADValues[2076*12 +: 12], 32, 28, comp929minVal, comp929minI, comp929minJ);
    wire [11:0] comp930minVal;
    wire [5:0] comp930minI, comp930minJ;
    Comparator comp930(SADValues[2013*12 +: 12], 31, 29, SADValues[1950*12 +: 12], 30, 30, comp930minVal, comp930minI, comp930minJ);
    wire [11:0] comp931minVal;
    wire [5:0] comp931minI, comp931minJ;
    Comparator comp931(SADValues[1887*12 +: 12], 29, 31, SADValues[1824*12 +: 12], 28, 32, comp931minVal, comp931minI, comp931minJ);
    wire [11:0] comp932minVal;
    wire [5:0] comp932minI, comp932minJ;
    Comparator comp932(SADValues[1761*12 +: 12], 27, 33, SADValues[1698*12 +: 12], 26, 34, comp932minVal, comp932minI, comp932minJ);
    wire [11:0] comp933minVal;
    wire [5:0] comp933minI, comp933minJ;
    Comparator comp933(SADValues[1635*12 +: 12], 25, 35, SADValues[1572*12 +: 12], 24, 36, comp933minVal, comp933minI, comp933minJ);
    wire [11:0] comp934minVal;
    wire [5:0] comp934minI, comp934minJ;
    Comparator comp934(SADValues[1509*12 +: 12], 23, 37, SADValues[1446*12 +: 12], 22, 38, comp934minVal, comp934minI, comp934minJ);
    wire [11:0] comp935minVal;
    wire [5:0] comp935minI, comp935minJ;
    Comparator comp935(SADValues[1383*12 +: 12], 21, 39, SADValues[1320*12 +: 12], 20, 40, comp935minVal, comp935minI, comp935minJ);
    wire [11:0] comp936minVal;
    wire [5:0] comp936minI, comp936minJ;
    Comparator comp936(SADValues[1257*12 +: 12], 19, 41, SADValues[1194*12 +: 12], 18, 42, comp936minVal, comp936minI, comp936minJ);
    wire [11:0] comp937minVal;
    wire [5:0] comp937minI, comp937minJ;
    Comparator comp937(SADValues[1131*12 +: 12], 17, 43, SADValues[1068*12 +: 12], 16, 44, comp937minVal, comp937minI, comp937minJ);
    wire [11:0] comp938minVal;
    wire [5:0] comp938minI, comp938minJ;
    Comparator comp938(SADValues[1005*12 +: 12], 15, 45, SADValues[942*12 +: 12], 14, 46, comp938minVal, comp938minI, comp938minJ);
    wire [11:0] comp939minVal;
    wire [5:0] comp939minI, comp939minJ;
    Comparator comp939(SADValues[879*12 +: 12], 13, 47, SADValues[816*12 +: 12], 12, 48, comp939minVal, comp939minI, comp939minJ);
    wire [11:0] comp940minVal;
    wire [5:0] comp940minI, comp940minJ;
    Comparator comp940(SADValues[753*12 +: 12], 11, 49, SADValues[690*12 +: 12], 10, 50, comp940minVal, comp940minI, comp940minJ);
    wire [11:0] comp941minVal;
    wire [5:0] comp941minI, comp941minJ;
    Comparator comp941(SADValues[627*12 +: 12], 9, 51, SADValues[564*12 +: 12], 8, 52, comp941minVal, comp941minI, comp941minJ);
    wire [11:0] comp942minVal;
    wire [5:0] comp942minI, comp942minJ;
    Comparator comp942(SADValues[501*12 +: 12], 7, 53, SADValues[438*12 +: 12], 6, 54, comp942minVal, comp942minI, comp942minJ);
    wire [11:0] comp943minVal;
    wire [5:0] comp943minI, comp943minJ;
    Comparator comp943(SADValues[375*12 +: 12], 5, 55, SADValues[312*12 +: 12], 4, 56, comp943minVal, comp943minI, comp943minJ);
    wire [11:0] comp944minVal;
    wire [5:0] comp944minI, comp944minJ;
    Comparator comp944(SADValues[249*12 +: 12], 3, 57, SADValues[186*12 +: 12], 2, 58, comp944minVal, comp944minI, comp944minJ);
    wire [11:0] comp945minVal;
    wire [5:0] comp945minI, comp945minJ;
    Comparator comp945(SADValues[123*12 +: 12], 1, 59, SADValues[60*12 +: 12], 0, 60, comp945minVal, comp945minI, comp945minJ);
    wire [11:0] comp946minVal;
    wire [5:0] comp946minI, comp946minJ;
    Comparator comp946(SADValues[124*12 +: 12], 1, 60, SADValues[187*12 +: 12], 2, 59, comp946minVal, comp946minI, comp946minJ);
    wire [11:0] comp947minVal;
    wire [5:0] comp947minI, comp947minJ;
    Comparator comp947(SADValues[250*12 +: 12], 3, 58, SADValues[313*12 +: 12], 4, 57, comp947minVal, comp947minI, comp947minJ);
    wire [11:0] comp948minVal;
    wire [5:0] comp948minI, comp948minJ;
    Comparator comp948(SADValues[376*12 +: 12], 5, 56, SADValues[439*12 +: 12], 6, 55, comp948minVal, comp948minI, comp948minJ);
    wire [11:0] comp949minVal;
    wire [5:0] comp949minI, comp949minJ;
    Comparator comp949(SADValues[502*12 +: 12], 7, 54, SADValues[565*12 +: 12], 8, 53, comp949minVal, comp949minI, comp949minJ);
    wire [11:0] comp950minVal;
    wire [5:0] comp950minI, comp950minJ;
    Comparator comp950(SADValues[628*12 +: 12], 9, 52, SADValues[691*12 +: 12], 10, 51, comp950minVal, comp950minI, comp950minJ);
    wire [11:0] comp951minVal;
    wire [5:0] comp951minI, comp951minJ;
    Comparator comp951(SADValues[754*12 +: 12], 11, 50, SADValues[817*12 +: 12], 12, 49, comp951minVal, comp951minI, comp951minJ);
    wire [11:0] comp952minVal;
    wire [5:0] comp952minI, comp952minJ;
    Comparator comp952(SADValues[880*12 +: 12], 13, 48, SADValues[943*12 +: 12], 14, 47, comp952minVal, comp952minI, comp952minJ);
    wire [11:0] comp953minVal;
    wire [5:0] comp953minI, comp953minJ;
    Comparator comp953(SADValues[1006*12 +: 12], 15, 46, SADValues[1069*12 +: 12], 16, 45, comp953minVal, comp953minI, comp953minJ);
    wire [11:0] comp954minVal;
    wire [5:0] comp954minI, comp954minJ;
    Comparator comp954(SADValues[1132*12 +: 12], 17, 44, SADValues[1195*12 +: 12], 18, 43, comp954minVal, comp954minI, comp954minJ);
    wire [11:0] comp955minVal;
    wire [5:0] comp955minI, comp955minJ;
    Comparator comp955(SADValues[1258*12 +: 12], 19, 42, SADValues[1321*12 +: 12], 20, 41, comp955minVal, comp955minI, comp955minJ);
    wire [11:0] comp956minVal;
    wire [5:0] comp956minI, comp956minJ;
    Comparator comp956(SADValues[1384*12 +: 12], 21, 40, SADValues[1447*12 +: 12], 22, 39, comp956minVal, comp956minI, comp956minJ);
    wire [11:0] comp957minVal;
    wire [5:0] comp957minI, comp957minJ;
    Comparator comp957(SADValues[1510*12 +: 12], 23, 38, SADValues[1573*12 +: 12], 24, 37, comp957minVal, comp957minI, comp957minJ);
    wire [11:0] comp958minVal;
    wire [5:0] comp958minI, comp958minJ;
    Comparator comp958(SADValues[1636*12 +: 12], 25, 36, SADValues[1699*12 +: 12], 26, 35, comp958minVal, comp958minI, comp958minJ);
    wire [11:0] comp959minVal;
    wire [5:0] comp959minI, comp959minJ;
    Comparator comp959(SADValues[1762*12 +: 12], 27, 34, SADValues[1825*12 +: 12], 28, 33, comp959minVal, comp959minI, comp959minJ);
    wire [11:0] comp960minVal;
    wire [5:0] comp960minI, comp960minJ;
    Comparator comp960(SADValues[1888*12 +: 12], 29, 32, SADValues[1951*12 +: 12], 30, 31, comp960minVal, comp960minI, comp960minJ);
    wire [11:0] comp961minVal;
    wire [5:0] comp961minI, comp961minJ;
    Comparator comp961(SADValues[2014*12 +: 12], 31, 30, SADValues[2077*12 +: 12], 32, 29, comp961minVal, comp961minI, comp961minJ);
    wire [11:0] comp962minVal;
    wire [5:0] comp962minI, comp962minJ;
    Comparator comp962(SADValues[2140*12 +: 12], 33, 28, SADValues[2203*12 +: 12], 34, 27, comp962minVal, comp962minI, comp962minJ);
    wire [11:0] comp963minVal;
    wire [5:0] comp963minI, comp963minJ;
    Comparator comp963(SADValues[2266*12 +: 12], 35, 26, SADValues[2329*12 +: 12], 36, 25, comp963minVal, comp963minI, comp963minJ);
    wire [11:0] comp964minVal;
    wire [5:0] comp964minI, comp964minJ;
    Comparator comp964(SADValues[2392*12 +: 12], 37, 24, SADValues[2455*12 +: 12], 38, 23, comp964minVal, comp964minI, comp964minJ);
    wire [11:0] comp965minVal;
    wire [5:0] comp965minI, comp965minJ;
    Comparator comp965(SADValues[2518*12 +: 12], 39, 22, SADValues[2581*12 +: 12], 40, 21, comp965minVal, comp965minI, comp965minJ);
    wire [11:0] comp966minVal;
    wire [5:0] comp966minI, comp966minJ;
    Comparator comp966(SADValues[2644*12 +: 12], 41, 20, SADValues[2707*12 +: 12], 42, 19, comp966minVal, comp966minI, comp966minJ);
    wire [11:0] comp967minVal;
    wire [5:0] comp967minI, comp967minJ;
    Comparator comp967(SADValues[2770*12 +: 12], 43, 18, SADValues[2833*12 +: 12], 44, 17, comp967minVal, comp967minI, comp967minJ);
    wire [11:0] comp968minVal;
    wire [5:0] comp968minI, comp968minJ;
    Comparator comp968(SADValues[2896*12 +: 12], 45, 16, SADValues[2959*12 +: 12], 46, 15, comp968minVal, comp968minI, comp968minJ);
    wire [11:0] comp969minVal;
    wire [5:0] comp969minI, comp969minJ;
    Comparator comp969(SADValues[3022*12 +: 12], 47, 14, SADValues[3085*12 +: 12], 48, 13, comp969minVal, comp969minI, comp969minJ);
    wire [11:0] comp970minVal;
    wire [5:0] comp970minI, comp970minJ;
    Comparator comp970(SADValues[3148*12 +: 12], 49, 12, SADValues[3211*12 +: 12], 50, 11, comp970minVal, comp970minI, comp970minJ);
    wire [11:0] comp971minVal;
    wire [5:0] comp971minI, comp971minJ;
    Comparator comp971(SADValues[3274*12 +: 12], 51, 10, SADValues[3337*12 +: 12], 52, 9, comp971minVal, comp971minI, comp971minJ);
    wire [11:0] comp972minVal;
    wire [5:0] comp972minI, comp972minJ;
    Comparator comp972(SADValues[3400*12 +: 12], 53, 8, SADValues[3463*12 +: 12], 54, 7, comp972minVal, comp972minI, comp972minJ);
    wire [11:0] comp973minVal;
    wire [5:0] comp973minI, comp973minJ;
    Comparator comp973(SADValues[3526*12 +: 12], 55, 6, SADValues[3589*12 +: 12], 56, 5, comp973minVal, comp973minI, comp973minJ);
    wire [11:0] comp974minVal;
    wire [5:0] comp974minI, comp974minJ;
    Comparator comp974(SADValues[3652*12 +: 12], 57, 4, SADValues[3715*12 +: 12], 58, 3, comp974minVal, comp974minI, comp974minJ);
    wire [11:0] comp975minVal;
    wire [5:0] comp975minI, comp975minJ;
    Comparator comp975(SADValues[3778*12 +: 12], 59, 2, SADValues[3841*12 +: 12], 60, 1, comp975minVal, comp975minI, comp975minJ);
    wire [11:0] comp976minVal;
    wire [5:0] comp976minI, comp976minJ;
    Comparator comp976(SADValues[3842*12 +: 12], 60, 2, SADValues[3779*12 +: 12], 59, 3, comp976minVal, comp976minI, comp976minJ);
    wire [11:0] comp977minVal;
    wire [5:0] comp977minI, comp977minJ;
    Comparator comp977(SADValues[3716*12 +: 12], 58, 4, SADValues[3653*12 +: 12], 57, 5, comp977minVal, comp977minI, comp977minJ);
    wire [11:0] comp978minVal;
    wire [5:0] comp978minI, comp978minJ;
    Comparator comp978(SADValues[3590*12 +: 12], 56, 6, SADValues[3527*12 +: 12], 55, 7, comp978minVal, comp978minI, comp978minJ);
    wire [11:0] comp979minVal;
    wire [5:0] comp979minI, comp979minJ;
    Comparator comp979(SADValues[3464*12 +: 12], 54, 8, SADValues[3401*12 +: 12], 53, 9, comp979minVal, comp979minI, comp979minJ);
    wire [11:0] comp980minVal;
    wire [5:0] comp980minI, comp980minJ;
    Comparator comp980(SADValues[3338*12 +: 12], 52, 10, SADValues[3275*12 +: 12], 51, 11, comp980minVal, comp980minI, comp980minJ);
    wire [11:0] comp981minVal;
    wire [5:0] comp981minI, comp981minJ;
    Comparator comp981(SADValues[3212*12 +: 12], 50, 12, SADValues[3149*12 +: 12], 49, 13, comp981minVal, comp981minI, comp981minJ);
    wire [11:0] comp982minVal;
    wire [5:0] comp982minI, comp982minJ;
    Comparator comp982(SADValues[3086*12 +: 12], 48, 14, SADValues[3023*12 +: 12], 47, 15, comp982minVal, comp982minI, comp982minJ);
    wire [11:0] comp983minVal;
    wire [5:0] comp983minI, comp983minJ;
    Comparator comp983(SADValues[2960*12 +: 12], 46, 16, SADValues[2897*12 +: 12], 45, 17, comp983minVal, comp983minI, comp983minJ);
    wire [11:0] comp984minVal;
    wire [5:0] comp984minI, comp984minJ;
    Comparator comp984(SADValues[2834*12 +: 12], 44, 18, SADValues[2771*12 +: 12], 43, 19, comp984minVal, comp984minI, comp984minJ);
    wire [11:0] comp985minVal;
    wire [5:0] comp985minI, comp985minJ;
    Comparator comp985(SADValues[2708*12 +: 12], 42, 20, SADValues[2645*12 +: 12], 41, 21, comp985minVal, comp985minI, comp985minJ);
    wire [11:0] comp986minVal;
    wire [5:0] comp986minI, comp986minJ;
    Comparator comp986(SADValues[2582*12 +: 12], 40, 22, SADValues[2519*12 +: 12], 39, 23, comp986minVal, comp986minI, comp986minJ);
    wire [11:0] comp987minVal;
    wire [5:0] comp987minI, comp987minJ;
    Comparator comp987(SADValues[2456*12 +: 12], 38, 24, SADValues[2393*12 +: 12], 37, 25, comp987minVal, comp987minI, comp987minJ);
    wire [11:0] comp988minVal;
    wire [5:0] comp988minI, comp988minJ;
    Comparator comp988(SADValues[2330*12 +: 12], 36, 26, SADValues[2267*12 +: 12], 35, 27, comp988minVal, comp988minI, comp988minJ);
    wire [11:0] comp989minVal;
    wire [5:0] comp989minI, comp989minJ;
    Comparator comp989(SADValues[2204*12 +: 12], 34, 28, SADValues[2141*12 +: 12], 33, 29, comp989minVal, comp989minI, comp989minJ);
    wire [11:0] comp990minVal;
    wire [5:0] comp990minI, comp990minJ;
    Comparator comp990(SADValues[2078*12 +: 12], 32, 30, SADValues[2015*12 +: 12], 31, 31, comp990minVal, comp990minI, comp990minJ);
    wire [11:0] comp991minVal;
    wire [5:0] comp991minI, comp991minJ;
    Comparator comp991(SADValues[1952*12 +: 12], 30, 32, SADValues[1889*12 +: 12], 29, 33, comp991minVal, comp991minI, comp991minJ);
    wire [11:0] comp992minVal;
    wire [5:0] comp992minI, comp992minJ;
    Comparator comp992(SADValues[1826*12 +: 12], 28, 34, SADValues[1763*12 +: 12], 27, 35, comp992minVal, comp992minI, comp992minJ);
    wire [11:0] comp993minVal;
    wire [5:0] comp993minI, comp993minJ;
    Comparator comp993(SADValues[1700*12 +: 12], 26, 36, SADValues[1637*12 +: 12], 25, 37, comp993minVal, comp993minI, comp993minJ);
    wire [11:0] comp994minVal;
    wire [5:0] comp994minI, comp994minJ;
    Comparator comp994(SADValues[1574*12 +: 12], 24, 38, SADValues[1511*12 +: 12], 23, 39, comp994minVal, comp994minI, comp994minJ);
    wire [11:0] comp995minVal;
    wire [5:0] comp995minI, comp995minJ;
    Comparator comp995(SADValues[1448*12 +: 12], 22, 40, SADValues[1385*12 +: 12], 21, 41, comp995minVal, comp995minI, comp995minJ);
    wire [11:0] comp996minVal;
    wire [5:0] comp996minI, comp996minJ;
    Comparator comp996(SADValues[1322*12 +: 12], 20, 42, SADValues[1259*12 +: 12], 19, 43, comp996minVal, comp996minI, comp996minJ);
    wire [11:0] comp997minVal;
    wire [5:0] comp997minI, comp997minJ;
    Comparator comp997(SADValues[1196*12 +: 12], 18, 44, SADValues[1133*12 +: 12], 17, 45, comp997minVal, comp997minI, comp997minJ);
    wire [11:0] comp998minVal;
    wire [5:0] comp998minI, comp998minJ;
    Comparator comp998(SADValues[1070*12 +: 12], 16, 46, SADValues[1007*12 +: 12], 15, 47, comp998minVal, comp998minI, comp998minJ);
    wire [11:0] comp999minVal;
    wire [5:0] comp999minI, comp999minJ;
    Comparator comp999(SADValues[944*12 +: 12], 14, 48, SADValues[881*12 +: 12], 13, 49, comp999minVal, comp999minI, comp999minJ);
    wire [11:0] comp1000minVal;
    wire [5:0] comp1000minI, comp1000minJ;
    Comparator comp1000(SADValues[818*12 +: 12], 12, 50, SADValues[755*12 +: 12], 11, 51, comp1000minVal, comp1000minI, comp1000minJ);
    wire [11:0] comp1001minVal;
    wire [5:0] comp1001minI, comp1001minJ;
    Comparator comp1001(SADValues[692*12 +: 12], 10, 52, SADValues[629*12 +: 12], 9, 53, comp1001minVal, comp1001minI, comp1001minJ);
    wire [11:0] comp1002minVal;
    wire [5:0] comp1002minI, comp1002minJ;
    Comparator comp1002(SADValues[566*12 +: 12], 8, 54, SADValues[503*12 +: 12], 7, 55, comp1002minVal, comp1002minI, comp1002minJ);
    wire [11:0] comp1003minVal;
    wire [5:0] comp1003minI, comp1003minJ;
    Comparator comp1003(SADValues[440*12 +: 12], 6, 56, SADValues[377*12 +: 12], 5, 57, comp1003minVal, comp1003minI, comp1003minJ);
    wire [11:0] comp1004minVal;
    wire [5:0] comp1004minI, comp1004minJ;
    Comparator comp1004(SADValues[314*12 +: 12], 4, 58, SADValues[251*12 +: 12], 3, 59, comp1004minVal, comp1004minI, comp1004minJ);
    wire [11:0] comp1005minVal;
    wire [5:0] comp1005minI, comp1005minJ;
    Comparator comp1005(SADValues[188*12 +: 12], 2, 60, SADValues[252*12 +: 12], 3, 60, comp1005minVal, comp1005minI, comp1005minJ);
    wire [11:0] comp1006minVal;
    wire [5:0] comp1006minI, comp1006minJ;
    Comparator comp1006(SADValues[315*12 +: 12], 4, 59, SADValues[378*12 +: 12], 5, 58, comp1006minVal, comp1006minI, comp1006minJ);
    wire [11:0] comp1007minVal;
    wire [5:0] comp1007minI, comp1007minJ;
    Comparator comp1007(SADValues[441*12 +: 12], 6, 57, SADValues[504*12 +: 12], 7, 56, comp1007minVal, comp1007minI, comp1007minJ);
    wire [11:0] comp1008minVal;
    wire [5:0] comp1008minI, comp1008minJ;
    Comparator comp1008(SADValues[567*12 +: 12], 8, 55, SADValues[630*12 +: 12], 9, 54, comp1008minVal, comp1008minI, comp1008minJ);
    wire [11:0] comp1009minVal;
    wire [5:0] comp1009minI, comp1009minJ;
    Comparator comp1009(SADValues[693*12 +: 12], 10, 53, SADValues[756*12 +: 12], 11, 52, comp1009minVal, comp1009minI, comp1009minJ);
    wire [11:0] comp1010minVal;
    wire [5:0] comp1010minI, comp1010minJ;
    Comparator comp1010(SADValues[819*12 +: 12], 12, 51, SADValues[882*12 +: 12], 13, 50, comp1010minVal, comp1010minI, comp1010minJ);
    wire [11:0] comp1011minVal;
    wire [5:0] comp1011minI, comp1011minJ;
    Comparator comp1011(SADValues[945*12 +: 12], 14, 49, SADValues[1008*12 +: 12], 15, 48, comp1011minVal, comp1011minI, comp1011minJ);
    wire [11:0] comp1012minVal;
    wire [5:0] comp1012minI, comp1012minJ;
    Comparator comp1012(SADValues[1071*12 +: 12], 16, 47, SADValues[1134*12 +: 12], 17, 46, comp1012minVal, comp1012minI, comp1012minJ);
    wire [11:0] comp1013minVal;
    wire [5:0] comp1013minI, comp1013minJ;
    Comparator comp1013(SADValues[1197*12 +: 12], 18, 45, SADValues[1260*12 +: 12], 19, 44, comp1013minVal, comp1013minI, comp1013minJ);
    wire [11:0] comp1014minVal;
    wire [5:0] comp1014minI, comp1014minJ;
    Comparator comp1014(SADValues[1323*12 +: 12], 20, 43, SADValues[1386*12 +: 12], 21, 42, comp1014minVal, comp1014minI, comp1014minJ);
    wire [11:0] comp1015minVal;
    wire [5:0] comp1015minI, comp1015minJ;
    Comparator comp1015(SADValues[1449*12 +: 12], 22, 41, SADValues[1512*12 +: 12], 23, 40, comp1015minVal, comp1015minI, comp1015minJ);
    wire [11:0] comp1016minVal;
    wire [5:0] comp1016minI, comp1016minJ;
    Comparator comp1016(SADValues[1575*12 +: 12], 24, 39, SADValues[1638*12 +: 12], 25, 38, comp1016minVal, comp1016minI, comp1016minJ);
    wire [11:0] comp1017minVal;
    wire [5:0] comp1017minI, comp1017minJ;
    Comparator comp1017(SADValues[1701*12 +: 12], 26, 37, SADValues[1764*12 +: 12], 27, 36, comp1017minVal, comp1017minI, comp1017minJ);
    wire [11:0] comp1018minVal;
    wire [5:0] comp1018minI, comp1018minJ;
    Comparator comp1018(SADValues[1827*12 +: 12], 28, 35, SADValues[1890*12 +: 12], 29, 34, comp1018minVal, comp1018minI, comp1018minJ);
    wire [11:0] comp1019minVal;
    wire [5:0] comp1019minI, comp1019minJ;
    Comparator comp1019(SADValues[1953*12 +: 12], 30, 33, SADValues[2016*12 +: 12], 31, 32, comp1019minVal, comp1019minI, comp1019minJ);
    wire [11:0] comp1020minVal;
    wire [5:0] comp1020minI, comp1020minJ;
    Comparator comp1020(SADValues[2079*12 +: 12], 32, 31, SADValues[2142*12 +: 12], 33, 30, comp1020minVal, comp1020minI, comp1020minJ);
    wire [11:0] comp1021minVal;
    wire [5:0] comp1021minI, comp1021minJ;
    Comparator comp1021(SADValues[2205*12 +: 12], 34, 29, SADValues[2268*12 +: 12], 35, 28, comp1021minVal, comp1021minI, comp1021minJ);
    wire [11:0] comp1022minVal;
    wire [5:0] comp1022minI, comp1022minJ;
    Comparator comp1022(SADValues[2331*12 +: 12], 36, 27, SADValues[2394*12 +: 12], 37, 26, comp1022minVal, comp1022minI, comp1022minJ);
    wire [11:0] comp1023minVal;
    wire [5:0] comp1023minI, comp1023minJ;
    Comparator comp1023(SADValues[2457*12 +: 12], 38, 25, SADValues[2520*12 +: 12], 39, 24, comp1023minVal, comp1023minI, comp1023minJ);
    wire [11:0] comp1024minVal;
    wire [5:0] comp1024minI, comp1024minJ;
    Comparator comp1024(SADValues[2583*12 +: 12], 40, 23, SADValues[2646*12 +: 12], 41, 22, comp1024minVal, comp1024minI, comp1024minJ);
    wire [11:0] comp1025minVal;
    wire [5:0] comp1025minI, comp1025minJ;
    Comparator comp1025(SADValues[2709*12 +: 12], 42, 21, SADValues[2772*12 +: 12], 43, 20, comp1025minVal, comp1025minI, comp1025minJ);
    wire [11:0] comp1026minVal;
    wire [5:0] comp1026minI, comp1026minJ;
    Comparator comp1026(SADValues[2835*12 +: 12], 44, 19, SADValues[2898*12 +: 12], 45, 18, comp1026minVal, comp1026minI, comp1026minJ);
    wire [11:0] comp1027minVal;
    wire [5:0] comp1027minI, comp1027minJ;
    Comparator comp1027(SADValues[2961*12 +: 12], 46, 17, SADValues[3024*12 +: 12], 47, 16, comp1027minVal, comp1027minI, comp1027minJ);
    wire [11:0] comp1028minVal;
    wire [5:0] comp1028minI, comp1028minJ;
    Comparator comp1028(SADValues[3087*12 +: 12], 48, 15, SADValues[3150*12 +: 12], 49, 14, comp1028minVal, comp1028minI, comp1028minJ);
    wire [11:0] comp1029minVal;
    wire [5:0] comp1029minI, comp1029minJ;
    Comparator comp1029(SADValues[3213*12 +: 12], 50, 13, SADValues[3276*12 +: 12], 51, 12, comp1029minVal, comp1029minI, comp1029minJ);
    wire [11:0] comp1030minVal;
    wire [5:0] comp1030minI, comp1030minJ;
    Comparator comp1030(SADValues[3339*12 +: 12], 52, 11, SADValues[3402*12 +: 12], 53, 10, comp1030minVal, comp1030minI, comp1030minJ);
    wire [11:0] comp1031minVal;
    wire [5:0] comp1031minI, comp1031minJ;
    Comparator comp1031(SADValues[3465*12 +: 12], 54, 9, SADValues[3528*12 +: 12], 55, 8, comp1031minVal, comp1031minI, comp1031minJ);
    wire [11:0] comp1032minVal;
    wire [5:0] comp1032minI, comp1032minJ;
    Comparator comp1032(SADValues[3591*12 +: 12], 56, 7, SADValues[3654*12 +: 12], 57, 6, comp1032minVal, comp1032minI, comp1032minJ);
    wire [11:0] comp1033minVal;
    wire [5:0] comp1033minI, comp1033minJ;
    Comparator comp1033(SADValues[3717*12 +: 12], 58, 5, SADValues[3780*12 +: 12], 59, 4, comp1033minVal, comp1033minI, comp1033minJ);
    wire [11:0] comp1034minVal;
    wire [5:0] comp1034minI, comp1034minJ;
    Comparator comp1034(SADValues[3843*12 +: 12], 60, 3, SADValues[3844*12 +: 12], 60, 4, comp1034minVal, comp1034minI, comp1034minJ);
    wire [11:0] comp1035minVal;
    wire [5:0] comp1035minI, comp1035minJ;
    Comparator comp1035(SADValues[3781*12 +: 12], 59, 5, SADValues[3718*12 +: 12], 58, 6, comp1035minVal, comp1035minI, comp1035minJ);
    wire [11:0] comp1036minVal;
    wire [5:0] comp1036minI, comp1036minJ;
    Comparator comp1036(SADValues[3655*12 +: 12], 57, 7, SADValues[3592*12 +: 12], 56, 8, comp1036minVal, comp1036minI, comp1036minJ);
    wire [11:0] comp1037minVal;
    wire [5:0] comp1037minI, comp1037minJ;
    Comparator comp1037(SADValues[3529*12 +: 12], 55, 9, SADValues[3466*12 +: 12], 54, 10, comp1037minVal, comp1037minI, comp1037minJ);
    wire [11:0] comp1038minVal;
    wire [5:0] comp1038minI, comp1038minJ;
    Comparator comp1038(SADValues[3403*12 +: 12], 53, 11, SADValues[3340*12 +: 12], 52, 12, comp1038minVal, comp1038minI, comp1038minJ);
    wire [11:0] comp1039minVal;
    wire [5:0] comp1039minI, comp1039minJ;
    Comparator comp1039(SADValues[3277*12 +: 12], 51, 13, SADValues[3214*12 +: 12], 50, 14, comp1039minVal, comp1039minI, comp1039minJ);
    wire [11:0] comp1040minVal;
    wire [5:0] comp1040minI, comp1040minJ;
    Comparator comp1040(SADValues[3151*12 +: 12], 49, 15, SADValues[3088*12 +: 12], 48, 16, comp1040minVal, comp1040minI, comp1040minJ);
    wire [11:0] comp1041minVal;
    wire [5:0] comp1041minI, comp1041minJ;
    Comparator comp1041(SADValues[3025*12 +: 12], 47, 17, SADValues[2962*12 +: 12], 46, 18, comp1041minVal, comp1041minI, comp1041minJ);
    wire [11:0] comp1042minVal;
    wire [5:0] comp1042minI, comp1042minJ;
    Comparator comp1042(SADValues[2899*12 +: 12], 45, 19, SADValues[2836*12 +: 12], 44, 20, comp1042minVal, comp1042minI, comp1042minJ);
    wire [11:0] comp1043minVal;
    wire [5:0] comp1043minI, comp1043minJ;
    Comparator comp1043(SADValues[2773*12 +: 12], 43, 21, SADValues[2710*12 +: 12], 42, 22, comp1043minVal, comp1043minI, comp1043minJ);
    wire [11:0] comp1044minVal;
    wire [5:0] comp1044minI, comp1044minJ;
    Comparator comp1044(SADValues[2647*12 +: 12], 41, 23, SADValues[2584*12 +: 12], 40, 24, comp1044minVal, comp1044minI, comp1044minJ);
    wire [11:0] comp1045minVal;
    wire [5:0] comp1045minI, comp1045minJ;
    Comparator comp1045(SADValues[2521*12 +: 12], 39, 25, SADValues[2458*12 +: 12], 38, 26, comp1045minVal, comp1045minI, comp1045minJ);
    wire [11:0] comp1046minVal;
    wire [5:0] comp1046minI, comp1046minJ;
    Comparator comp1046(SADValues[2395*12 +: 12], 37, 27, SADValues[2332*12 +: 12], 36, 28, comp1046minVal, comp1046minI, comp1046minJ);
    wire [11:0] comp1047minVal;
    wire [5:0] comp1047minI, comp1047minJ;
    Comparator comp1047(SADValues[2269*12 +: 12], 35, 29, SADValues[2206*12 +: 12], 34, 30, comp1047minVal, comp1047minI, comp1047minJ);
    wire [11:0] comp1048minVal;
    wire [5:0] comp1048minI, comp1048minJ;
    Comparator comp1048(SADValues[2143*12 +: 12], 33, 31, SADValues[2080*12 +: 12], 32, 32, comp1048minVal, comp1048minI, comp1048minJ);
    wire [11:0] comp1049minVal;
    wire [5:0] comp1049minI, comp1049minJ;
    Comparator comp1049(SADValues[2017*12 +: 12], 31, 33, SADValues[1954*12 +: 12], 30, 34, comp1049minVal, comp1049minI, comp1049minJ);
    wire [11:0] comp1050minVal;
    wire [5:0] comp1050minI, comp1050minJ;
    Comparator comp1050(SADValues[1891*12 +: 12], 29, 35, SADValues[1828*12 +: 12], 28, 36, comp1050minVal, comp1050minI, comp1050minJ);
    wire [11:0] comp1051minVal;
    wire [5:0] comp1051minI, comp1051minJ;
    Comparator comp1051(SADValues[1765*12 +: 12], 27, 37, SADValues[1702*12 +: 12], 26, 38, comp1051minVal, comp1051minI, comp1051minJ);
    wire [11:0] comp1052minVal;
    wire [5:0] comp1052minI, comp1052minJ;
    Comparator comp1052(SADValues[1639*12 +: 12], 25, 39, SADValues[1576*12 +: 12], 24, 40, comp1052minVal, comp1052minI, comp1052minJ);
    wire [11:0] comp1053minVal;
    wire [5:0] comp1053minI, comp1053minJ;
    Comparator comp1053(SADValues[1513*12 +: 12], 23, 41, SADValues[1450*12 +: 12], 22, 42, comp1053minVal, comp1053minI, comp1053minJ);
    wire [11:0] comp1054minVal;
    wire [5:0] comp1054minI, comp1054minJ;
    Comparator comp1054(SADValues[1387*12 +: 12], 21, 43, SADValues[1324*12 +: 12], 20, 44, comp1054minVal, comp1054minI, comp1054minJ);
    wire [11:0] comp1055minVal;
    wire [5:0] comp1055minI, comp1055minJ;
    Comparator comp1055(SADValues[1261*12 +: 12], 19, 45, SADValues[1198*12 +: 12], 18, 46, comp1055minVal, comp1055minI, comp1055minJ);
    wire [11:0] comp1056minVal;
    wire [5:0] comp1056minI, comp1056minJ;
    Comparator comp1056(SADValues[1135*12 +: 12], 17, 47, SADValues[1072*12 +: 12], 16, 48, comp1056minVal, comp1056minI, comp1056minJ);
    wire [11:0] comp1057minVal;
    wire [5:0] comp1057minI, comp1057minJ;
    Comparator comp1057(SADValues[1009*12 +: 12], 15, 49, SADValues[946*12 +: 12], 14, 50, comp1057minVal, comp1057minI, comp1057minJ);
    wire [11:0] comp1058minVal;
    wire [5:0] comp1058minI, comp1058minJ;
    Comparator comp1058(SADValues[883*12 +: 12], 13, 51, SADValues[820*12 +: 12], 12, 52, comp1058minVal, comp1058minI, comp1058minJ);
    wire [11:0] comp1059minVal;
    wire [5:0] comp1059minI, comp1059minJ;
    Comparator comp1059(SADValues[757*12 +: 12], 11, 53, SADValues[694*12 +: 12], 10, 54, comp1059minVal, comp1059minI, comp1059minJ);
    wire [11:0] comp1060minVal;
    wire [5:0] comp1060minI, comp1060minJ;
    Comparator comp1060(SADValues[631*12 +: 12], 9, 55, SADValues[568*12 +: 12], 8, 56, comp1060minVal, comp1060minI, comp1060minJ);
    wire [11:0] comp1061minVal;
    wire [5:0] comp1061minI, comp1061minJ;
    Comparator comp1061(SADValues[505*12 +: 12], 7, 57, SADValues[442*12 +: 12], 6, 58, comp1061minVal, comp1061minI, comp1061minJ);
    wire [11:0] comp1062minVal;
    wire [5:0] comp1062minI, comp1062minJ;
    Comparator comp1062(SADValues[379*12 +: 12], 5, 59, SADValues[316*12 +: 12], 4, 60, comp1062minVal, comp1062minI, comp1062minJ);
    wire [11:0] comp1063minVal;
    wire [5:0] comp1063minI, comp1063minJ;
    Comparator comp1063(SADValues[380*12 +: 12], 5, 60, SADValues[443*12 +: 12], 6, 59, comp1063minVal, comp1063minI, comp1063minJ);
    wire [11:0] comp1064minVal;
    wire [5:0] comp1064minI, comp1064minJ;
    Comparator comp1064(SADValues[506*12 +: 12], 7, 58, SADValues[569*12 +: 12], 8, 57, comp1064minVal, comp1064minI, comp1064minJ);
    wire [11:0] comp1065minVal;
    wire [5:0] comp1065minI, comp1065minJ;
    Comparator comp1065(SADValues[632*12 +: 12], 9, 56, SADValues[695*12 +: 12], 10, 55, comp1065minVal, comp1065minI, comp1065minJ);
    wire [11:0] comp1066minVal;
    wire [5:0] comp1066minI, comp1066minJ;
    Comparator comp1066(SADValues[758*12 +: 12], 11, 54, SADValues[821*12 +: 12], 12, 53, comp1066minVal, comp1066minI, comp1066minJ);
    wire [11:0] comp1067minVal;
    wire [5:0] comp1067minI, comp1067minJ;
    Comparator comp1067(SADValues[884*12 +: 12], 13, 52, SADValues[947*12 +: 12], 14, 51, comp1067minVal, comp1067minI, comp1067minJ);
    wire [11:0] comp1068minVal;
    wire [5:0] comp1068minI, comp1068minJ;
    Comparator comp1068(SADValues[1010*12 +: 12], 15, 50, SADValues[1073*12 +: 12], 16, 49, comp1068minVal, comp1068minI, comp1068minJ);
    wire [11:0] comp1069minVal;
    wire [5:0] comp1069minI, comp1069minJ;
    Comparator comp1069(SADValues[1136*12 +: 12], 17, 48, SADValues[1199*12 +: 12], 18, 47, comp1069minVal, comp1069minI, comp1069minJ);
    wire [11:0] comp1070minVal;
    wire [5:0] comp1070minI, comp1070minJ;
    Comparator comp1070(SADValues[1262*12 +: 12], 19, 46, SADValues[1325*12 +: 12], 20, 45, comp1070minVal, comp1070minI, comp1070minJ);
    wire [11:0] comp1071minVal;
    wire [5:0] comp1071minI, comp1071minJ;
    Comparator comp1071(SADValues[1388*12 +: 12], 21, 44, SADValues[1451*12 +: 12], 22, 43, comp1071minVal, comp1071minI, comp1071minJ);
    wire [11:0] comp1072minVal;
    wire [5:0] comp1072minI, comp1072minJ;
    Comparator comp1072(SADValues[1514*12 +: 12], 23, 42, SADValues[1577*12 +: 12], 24, 41, comp1072minVal, comp1072minI, comp1072minJ);
    wire [11:0] comp1073minVal;
    wire [5:0] comp1073minI, comp1073minJ;
    Comparator comp1073(SADValues[1640*12 +: 12], 25, 40, SADValues[1703*12 +: 12], 26, 39, comp1073minVal, comp1073minI, comp1073minJ);
    wire [11:0] comp1074minVal;
    wire [5:0] comp1074minI, comp1074minJ;
    Comparator comp1074(SADValues[1766*12 +: 12], 27, 38, SADValues[1829*12 +: 12], 28, 37, comp1074minVal, comp1074minI, comp1074minJ);
    wire [11:0] comp1075minVal;
    wire [5:0] comp1075minI, comp1075minJ;
    Comparator comp1075(SADValues[1892*12 +: 12], 29, 36, SADValues[1955*12 +: 12], 30, 35, comp1075minVal, comp1075minI, comp1075minJ);
    wire [11:0] comp1076minVal;
    wire [5:0] comp1076minI, comp1076minJ;
    Comparator comp1076(SADValues[2018*12 +: 12], 31, 34, SADValues[2081*12 +: 12], 32, 33, comp1076minVal, comp1076minI, comp1076minJ);
    wire [11:0] comp1077minVal;
    wire [5:0] comp1077minI, comp1077minJ;
    Comparator comp1077(SADValues[2144*12 +: 12], 33, 32, SADValues[2207*12 +: 12], 34, 31, comp1077minVal, comp1077minI, comp1077minJ);
    wire [11:0] comp1078minVal;
    wire [5:0] comp1078minI, comp1078minJ;
    Comparator comp1078(SADValues[2270*12 +: 12], 35, 30, SADValues[2333*12 +: 12], 36, 29, comp1078minVal, comp1078minI, comp1078minJ);
    wire [11:0] comp1079minVal;
    wire [5:0] comp1079minI, comp1079minJ;
    Comparator comp1079(SADValues[2396*12 +: 12], 37, 28, SADValues[2459*12 +: 12], 38, 27, comp1079minVal, comp1079minI, comp1079minJ);
    wire [11:0] comp1080minVal;
    wire [5:0] comp1080minI, comp1080minJ;
    Comparator comp1080(SADValues[2522*12 +: 12], 39, 26, SADValues[2585*12 +: 12], 40, 25, comp1080minVal, comp1080minI, comp1080minJ);
    wire [11:0] comp1081minVal;
    wire [5:0] comp1081minI, comp1081minJ;
    Comparator comp1081(SADValues[2648*12 +: 12], 41, 24, SADValues[2711*12 +: 12], 42, 23, comp1081minVal, comp1081minI, comp1081minJ);
    wire [11:0] comp1082minVal;
    wire [5:0] comp1082minI, comp1082minJ;
    Comparator comp1082(SADValues[2774*12 +: 12], 43, 22, SADValues[2837*12 +: 12], 44, 21, comp1082minVal, comp1082minI, comp1082minJ);
    wire [11:0] comp1083minVal;
    wire [5:0] comp1083minI, comp1083minJ;
    Comparator comp1083(SADValues[2900*12 +: 12], 45, 20, SADValues[2963*12 +: 12], 46, 19, comp1083minVal, comp1083minI, comp1083minJ);
    wire [11:0] comp1084minVal;
    wire [5:0] comp1084minI, comp1084minJ;
    Comparator comp1084(SADValues[3026*12 +: 12], 47, 18, SADValues[3089*12 +: 12], 48, 17, comp1084minVal, comp1084minI, comp1084minJ);
    wire [11:0] comp1085minVal;
    wire [5:0] comp1085minI, comp1085minJ;
    Comparator comp1085(SADValues[3152*12 +: 12], 49, 16, SADValues[3215*12 +: 12], 50, 15, comp1085minVal, comp1085minI, comp1085minJ);
    wire [11:0] comp1086minVal;
    wire [5:0] comp1086minI, comp1086minJ;
    Comparator comp1086(SADValues[3278*12 +: 12], 51, 14, SADValues[3341*12 +: 12], 52, 13, comp1086minVal, comp1086minI, comp1086minJ);
    wire [11:0] comp1087minVal;
    wire [5:0] comp1087minI, comp1087minJ;
    Comparator comp1087(SADValues[3404*12 +: 12], 53, 12, SADValues[3467*12 +: 12], 54, 11, comp1087minVal, comp1087minI, comp1087minJ);
    wire [11:0] comp1088minVal;
    wire [5:0] comp1088minI, comp1088minJ;
    Comparator comp1088(SADValues[3530*12 +: 12], 55, 10, SADValues[3593*12 +: 12], 56, 9, comp1088minVal, comp1088minI, comp1088minJ);
    wire [11:0] comp1089minVal;
    wire [5:0] comp1089minI, comp1089minJ;
    Comparator comp1089(SADValues[3656*12 +: 12], 57, 8, SADValues[3719*12 +: 12], 58, 7, comp1089minVal, comp1089minI, comp1089minJ);
    wire [11:0] comp1090minVal;
    wire [5:0] comp1090minI, comp1090minJ;
    Comparator comp1090(SADValues[3782*12 +: 12], 59, 6, SADValues[3845*12 +: 12], 60, 5, comp1090minVal, comp1090minI, comp1090minJ);
    wire [11:0] comp1091minVal;
    wire [5:0] comp1091minI, comp1091minJ;
    Comparator comp1091(SADValues[3846*12 +: 12], 60, 6, SADValues[3783*12 +: 12], 59, 7, comp1091minVal, comp1091minI, comp1091minJ);
    wire [11:0] comp1092minVal;
    wire [5:0] comp1092minI, comp1092minJ;
    Comparator comp1092(SADValues[3720*12 +: 12], 58, 8, SADValues[3657*12 +: 12], 57, 9, comp1092minVal, comp1092minI, comp1092minJ);
    wire [11:0] comp1093minVal;
    wire [5:0] comp1093minI, comp1093minJ;
    Comparator comp1093(SADValues[3594*12 +: 12], 56, 10, SADValues[3531*12 +: 12], 55, 11, comp1093minVal, comp1093minI, comp1093minJ);
    wire [11:0] comp1094minVal;
    wire [5:0] comp1094minI, comp1094minJ;
    Comparator comp1094(SADValues[3468*12 +: 12], 54, 12, SADValues[3405*12 +: 12], 53, 13, comp1094minVal, comp1094minI, comp1094minJ);
    wire [11:0] comp1095minVal;
    wire [5:0] comp1095minI, comp1095minJ;
    Comparator comp1095(SADValues[3342*12 +: 12], 52, 14, SADValues[3279*12 +: 12], 51, 15, comp1095minVal, comp1095minI, comp1095minJ);
    wire [11:0] comp1096minVal;
    wire [5:0] comp1096minI, comp1096minJ;
    Comparator comp1096(SADValues[3216*12 +: 12], 50, 16, SADValues[3153*12 +: 12], 49, 17, comp1096minVal, comp1096minI, comp1096minJ);
    wire [11:0] comp1097minVal;
    wire [5:0] comp1097minI, comp1097minJ;
    Comparator comp1097(SADValues[3090*12 +: 12], 48, 18, SADValues[3027*12 +: 12], 47, 19, comp1097minVal, comp1097minI, comp1097minJ);
    wire [11:0] comp1098minVal;
    wire [5:0] comp1098minI, comp1098minJ;
    Comparator comp1098(SADValues[2964*12 +: 12], 46, 20, SADValues[2901*12 +: 12], 45, 21, comp1098minVal, comp1098minI, comp1098minJ);
    wire [11:0] comp1099minVal;
    wire [5:0] comp1099minI, comp1099minJ;
    Comparator comp1099(SADValues[2838*12 +: 12], 44, 22, SADValues[2775*12 +: 12], 43, 23, comp1099minVal, comp1099minI, comp1099minJ);
    wire [11:0] comp1100minVal;
    wire [5:0] comp1100minI, comp1100minJ;
    Comparator comp1100(SADValues[2712*12 +: 12], 42, 24, SADValues[2649*12 +: 12], 41, 25, comp1100minVal, comp1100minI, comp1100minJ);
    wire [11:0] comp1101minVal;
    wire [5:0] comp1101minI, comp1101minJ;
    Comparator comp1101(SADValues[2586*12 +: 12], 40, 26, SADValues[2523*12 +: 12], 39, 27, comp1101minVal, comp1101minI, comp1101minJ);
    wire [11:0] comp1102minVal;
    wire [5:0] comp1102minI, comp1102minJ;
    Comparator comp1102(SADValues[2460*12 +: 12], 38, 28, SADValues[2397*12 +: 12], 37, 29, comp1102minVal, comp1102minI, comp1102minJ);
    wire [11:0] comp1103minVal;
    wire [5:0] comp1103minI, comp1103minJ;
    Comparator comp1103(SADValues[2334*12 +: 12], 36, 30, SADValues[2271*12 +: 12], 35, 31, comp1103minVal, comp1103minI, comp1103minJ);
    wire [11:0] comp1104minVal;
    wire [5:0] comp1104minI, comp1104minJ;
    Comparator comp1104(SADValues[2208*12 +: 12], 34, 32, SADValues[2145*12 +: 12], 33, 33, comp1104minVal, comp1104minI, comp1104minJ);
    wire [11:0] comp1105minVal;
    wire [5:0] comp1105minI, comp1105minJ;
    Comparator comp1105(SADValues[2082*12 +: 12], 32, 34, SADValues[2019*12 +: 12], 31, 35, comp1105minVal, comp1105minI, comp1105minJ);
    wire [11:0] comp1106minVal;
    wire [5:0] comp1106minI, comp1106minJ;
    Comparator comp1106(SADValues[1956*12 +: 12], 30, 36, SADValues[1893*12 +: 12], 29, 37, comp1106minVal, comp1106minI, comp1106minJ);
    wire [11:0] comp1107minVal;
    wire [5:0] comp1107minI, comp1107minJ;
    Comparator comp1107(SADValues[1830*12 +: 12], 28, 38, SADValues[1767*12 +: 12], 27, 39, comp1107minVal, comp1107minI, comp1107minJ);
    wire [11:0] comp1108minVal;
    wire [5:0] comp1108minI, comp1108minJ;
    Comparator comp1108(SADValues[1704*12 +: 12], 26, 40, SADValues[1641*12 +: 12], 25, 41, comp1108minVal, comp1108minI, comp1108minJ);
    wire [11:0] comp1109minVal;
    wire [5:0] comp1109minI, comp1109minJ;
    Comparator comp1109(SADValues[1578*12 +: 12], 24, 42, SADValues[1515*12 +: 12], 23, 43, comp1109minVal, comp1109minI, comp1109minJ);
    wire [11:0] comp1110minVal;
    wire [5:0] comp1110minI, comp1110minJ;
    Comparator comp1110(SADValues[1452*12 +: 12], 22, 44, SADValues[1389*12 +: 12], 21, 45, comp1110minVal, comp1110minI, comp1110minJ);
    wire [11:0] comp1111minVal;
    wire [5:0] comp1111minI, comp1111minJ;
    Comparator comp1111(SADValues[1326*12 +: 12], 20, 46, SADValues[1263*12 +: 12], 19, 47, comp1111minVal, comp1111minI, comp1111minJ);
    wire [11:0] comp1112minVal;
    wire [5:0] comp1112minI, comp1112minJ;
    Comparator comp1112(SADValues[1200*12 +: 12], 18, 48, SADValues[1137*12 +: 12], 17, 49, comp1112minVal, comp1112minI, comp1112minJ);
    wire [11:0] comp1113minVal;
    wire [5:0] comp1113minI, comp1113minJ;
    Comparator comp1113(SADValues[1074*12 +: 12], 16, 50, SADValues[1011*12 +: 12], 15, 51, comp1113minVal, comp1113minI, comp1113minJ);
    wire [11:0] comp1114minVal;
    wire [5:0] comp1114minI, comp1114minJ;
    Comparator comp1114(SADValues[948*12 +: 12], 14, 52, SADValues[885*12 +: 12], 13, 53, comp1114minVal, comp1114minI, comp1114minJ);
    wire [11:0] comp1115minVal;
    wire [5:0] comp1115minI, comp1115minJ;
    Comparator comp1115(SADValues[822*12 +: 12], 12, 54, SADValues[759*12 +: 12], 11, 55, comp1115minVal, comp1115minI, comp1115minJ);
    wire [11:0] comp1116minVal;
    wire [5:0] comp1116minI, comp1116minJ;
    Comparator comp1116(SADValues[696*12 +: 12], 10, 56, SADValues[633*12 +: 12], 9, 57, comp1116minVal, comp1116minI, comp1116minJ);
    wire [11:0] comp1117minVal;
    wire [5:0] comp1117minI, comp1117minJ;
    Comparator comp1117(SADValues[570*12 +: 12], 8, 58, SADValues[507*12 +: 12], 7, 59, comp1117minVal, comp1117minI, comp1117minJ);
    wire [11:0] comp1118minVal;
    wire [5:0] comp1118minI, comp1118minJ;
    Comparator comp1118(SADValues[444*12 +: 12], 6, 60, SADValues[508*12 +: 12], 7, 60, comp1118minVal, comp1118minI, comp1118minJ);
    wire [11:0] comp1119minVal;
    wire [5:0] comp1119minI, comp1119minJ;
    Comparator comp1119(SADValues[571*12 +: 12], 8, 59, SADValues[634*12 +: 12], 9, 58, comp1119minVal, comp1119minI, comp1119minJ);
    wire [11:0] comp1120minVal;
    wire [5:0] comp1120minI, comp1120minJ;
    Comparator comp1120(SADValues[697*12 +: 12], 10, 57, SADValues[760*12 +: 12], 11, 56, comp1120minVal, comp1120minI, comp1120minJ);
    wire [11:0] comp1121minVal;
    wire [5:0] comp1121minI, comp1121minJ;
    Comparator comp1121(SADValues[823*12 +: 12], 12, 55, SADValues[886*12 +: 12], 13, 54, comp1121minVal, comp1121minI, comp1121minJ);
    wire [11:0] comp1122minVal;
    wire [5:0] comp1122minI, comp1122minJ;
    Comparator comp1122(SADValues[949*12 +: 12], 14, 53, SADValues[1012*12 +: 12], 15, 52, comp1122minVal, comp1122minI, comp1122minJ);
    wire [11:0] comp1123minVal;
    wire [5:0] comp1123minI, comp1123minJ;
    Comparator comp1123(SADValues[1075*12 +: 12], 16, 51, SADValues[1138*12 +: 12], 17, 50, comp1123minVal, comp1123minI, comp1123minJ);
    wire [11:0] comp1124minVal;
    wire [5:0] comp1124minI, comp1124minJ;
    Comparator comp1124(SADValues[1201*12 +: 12], 18, 49, SADValues[1264*12 +: 12], 19, 48, comp1124minVal, comp1124minI, comp1124minJ);
    wire [11:0] comp1125minVal;
    wire [5:0] comp1125minI, comp1125minJ;
    Comparator comp1125(SADValues[1327*12 +: 12], 20, 47, SADValues[1390*12 +: 12], 21, 46, comp1125minVal, comp1125minI, comp1125minJ);
    wire [11:0] comp1126minVal;
    wire [5:0] comp1126minI, comp1126minJ;
    Comparator comp1126(SADValues[1453*12 +: 12], 22, 45, SADValues[1516*12 +: 12], 23, 44, comp1126minVal, comp1126minI, comp1126minJ);
    wire [11:0] comp1127minVal;
    wire [5:0] comp1127minI, comp1127minJ;
    Comparator comp1127(SADValues[1579*12 +: 12], 24, 43, SADValues[1642*12 +: 12], 25, 42, comp1127minVal, comp1127minI, comp1127minJ);
    wire [11:0] comp1128minVal;
    wire [5:0] comp1128minI, comp1128minJ;
    Comparator comp1128(SADValues[1705*12 +: 12], 26, 41, SADValues[1768*12 +: 12], 27, 40, comp1128minVal, comp1128minI, comp1128minJ);
    wire [11:0] comp1129minVal;
    wire [5:0] comp1129minI, comp1129minJ;
    Comparator comp1129(SADValues[1831*12 +: 12], 28, 39, SADValues[1894*12 +: 12], 29, 38, comp1129minVal, comp1129minI, comp1129minJ);
    wire [11:0] comp1130minVal;
    wire [5:0] comp1130minI, comp1130minJ;
    Comparator comp1130(SADValues[1957*12 +: 12], 30, 37, SADValues[2020*12 +: 12], 31, 36, comp1130minVal, comp1130minI, comp1130minJ);
    wire [11:0] comp1131minVal;
    wire [5:0] comp1131minI, comp1131minJ;
    Comparator comp1131(SADValues[2083*12 +: 12], 32, 35, SADValues[2146*12 +: 12], 33, 34, comp1131minVal, comp1131minI, comp1131minJ);
    wire [11:0] comp1132minVal;
    wire [5:0] comp1132minI, comp1132minJ;
    Comparator comp1132(SADValues[2209*12 +: 12], 34, 33, SADValues[2272*12 +: 12], 35, 32, comp1132minVal, comp1132minI, comp1132minJ);
    wire [11:0] comp1133minVal;
    wire [5:0] comp1133minI, comp1133minJ;
    Comparator comp1133(SADValues[2335*12 +: 12], 36, 31, SADValues[2398*12 +: 12], 37, 30, comp1133minVal, comp1133minI, comp1133minJ);
    wire [11:0] comp1134minVal;
    wire [5:0] comp1134minI, comp1134minJ;
    Comparator comp1134(SADValues[2461*12 +: 12], 38, 29, SADValues[2524*12 +: 12], 39, 28, comp1134minVal, comp1134minI, comp1134minJ);
    wire [11:0] comp1135minVal;
    wire [5:0] comp1135minI, comp1135minJ;
    Comparator comp1135(SADValues[2587*12 +: 12], 40, 27, SADValues[2650*12 +: 12], 41, 26, comp1135minVal, comp1135minI, comp1135minJ);
    wire [11:0] comp1136minVal;
    wire [5:0] comp1136minI, comp1136minJ;
    Comparator comp1136(SADValues[2713*12 +: 12], 42, 25, SADValues[2776*12 +: 12], 43, 24, comp1136minVal, comp1136minI, comp1136minJ);
    wire [11:0] comp1137minVal;
    wire [5:0] comp1137minI, comp1137minJ;
    Comparator comp1137(SADValues[2839*12 +: 12], 44, 23, SADValues[2902*12 +: 12], 45, 22, comp1137minVal, comp1137minI, comp1137minJ);
    wire [11:0] comp1138minVal;
    wire [5:0] comp1138minI, comp1138minJ;
    Comparator comp1138(SADValues[2965*12 +: 12], 46, 21, SADValues[3028*12 +: 12], 47, 20, comp1138minVal, comp1138minI, comp1138minJ);
    wire [11:0] comp1139minVal;
    wire [5:0] comp1139minI, comp1139minJ;
    Comparator comp1139(SADValues[3091*12 +: 12], 48, 19, SADValues[3154*12 +: 12], 49, 18, comp1139minVal, comp1139minI, comp1139minJ);
    wire [11:0] comp1140minVal;
    wire [5:0] comp1140minI, comp1140minJ;
    Comparator comp1140(SADValues[3217*12 +: 12], 50, 17, SADValues[3280*12 +: 12], 51, 16, comp1140minVal, comp1140minI, comp1140minJ);
    wire [11:0] comp1141minVal;
    wire [5:0] comp1141minI, comp1141minJ;
    Comparator comp1141(SADValues[3343*12 +: 12], 52, 15, SADValues[3406*12 +: 12], 53, 14, comp1141minVal, comp1141minI, comp1141minJ);
    wire [11:0] comp1142minVal;
    wire [5:0] comp1142minI, comp1142minJ;
    Comparator comp1142(SADValues[3469*12 +: 12], 54, 13, SADValues[3532*12 +: 12], 55, 12, comp1142minVal, comp1142minI, comp1142minJ);
    wire [11:0] comp1143minVal;
    wire [5:0] comp1143minI, comp1143minJ;
    Comparator comp1143(SADValues[3595*12 +: 12], 56, 11, SADValues[3658*12 +: 12], 57, 10, comp1143minVal, comp1143minI, comp1143minJ);
    wire [11:0] comp1144minVal;
    wire [5:0] comp1144minI, comp1144minJ;
    Comparator comp1144(SADValues[3721*12 +: 12], 58, 9, SADValues[3784*12 +: 12], 59, 8, comp1144minVal, comp1144minI, comp1144minJ);
    wire [11:0] comp1145minVal;
    wire [5:0] comp1145minI, comp1145minJ;
    Comparator comp1145(SADValues[3847*12 +: 12], 60, 7, SADValues[3848*12 +: 12], 60, 8, comp1145minVal, comp1145minI, comp1145minJ);
    wire [11:0] comp1146minVal;
    wire [5:0] comp1146minI, comp1146minJ;
    Comparator comp1146(SADValues[3785*12 +: 12], 59, 9, SADValues[3722*12 +: 12], 58, 10, comp1146minVal, comp1146minI, comp1146minJ);
    wire [11:0] comp1147minVal;
    wire [5:0] comp1147minI, comp1147minJ;
    Comparator comp1147(SADValues[3659*12 +: 12], 57, 11, SADValues[3596*12 +: 12], 56, 12, comp1147minVal, comp1147minI, comp1147minJ);
    wire [11:0] comp1148minVal;
    wire [5:0] comp1148minI, comp1148minJ;
    Comparator comp1148(SADValues[3533*12 +: 12], 55, 13, SADValues[3470*12 +: 12], 54, 14, comp1148minVal, comp1148minI, comp1148minJ);
    wire [11:0] comp1149minVal;
    wire [5:0] comp1149minI, comp1149minJ;
    Comparator comp1149(SADValues[3407*12 +: 12], 53, 15, SADValues[3344*12 +: 12], 52, 16, comp1149minVal, comp1149minI, comp1149minJ);
    wire [11:0] comp1150minVal;
    wire [5:0] comp1150minI, comp1150minJ;
    Comparator comp1150(SADValues[3281*12 +: 12], 51, 17, SADValues[3218*12 +: 12], 50, 18, comp1150minVal, comp1150minI, comp1150minJ);
    wire [11:0] comp1151minVal;
    wire [5:0] comp1151minI, comp1151minJ;
    Comparator comp1151(SADValues[3155*12 +: 12], 49, 19, SADValues[3092*12 +: 12], 48, 20, comp1151minVal, comp1151minI, comp1151minJ);
    wire [11:0] comp1152minVal;
    wire [5:0] comp1152minI, comp1152minJ;
    Comparator comp1152(SADValues[3029*12 +: 12], 47, 21, SADValues[2966*12 +: 12], 46, 22, comp1152minVal, comp1152minI, comp1152minJ);
    wire [11:0] comp1153minVal;
    wire [5:0] comp1153minI, comp1153minJ;
    Comparator comp1153(SADValues[2903*12 +: 12], 45, 23, SADValues[2840*12 +: 12], 44, 24, comp1153minVal, comp1153minI, comp1153minJ);
    wire [11:0] comp1154minVal;
    wire [5:0] comp1154minI, comp1154minJ;
    Comparator comp1154(SADValues[2777*12 +: 12], 43, 25, SADValues[2714*12 +: 12], 42, 26, comp1154minVal, comp1154minI, comp1154minJ);
    wire [11:0] comp1155minVal;
    wire [5:0] comp1155minI, comp1155minJ;
    Comparator comp1155(SADValues[2651*12 +: 12], 41, 27, SADValues[2588*12 +: 12], 40, 28, comp1155minVal, comp1155minI, comp1155minJ);
    wire [11:0] comp1156minVal;
    wire [5:0] comp1156minI, comp1156minJ;
    Comparator comp1156(SADValues[2525*12 +: 12], 39, 29, SADValues[2462*12 +: 12], 38, 30, comp1156minVal, comp1156minI, comp1156minJ);
    wire [11:0] comp1157minVal;
    wire [5:0] comp1157minI, comp1157minJ;
    Comparator comp1157(SADValues[2399*12 +: 12], 37, 31, SADValues[2336*12 +: 12], 36, 32, comp1157minVal, comp1157minI, comp1157minJ);
    wire [11:0] comp1158minVal;
    wire [5:0] comp1158minI, comp1158minJ;
    Comparator comp1158(SADValues[2273*12 +: 12], 35, 33, SADValues[2210*12 +: 12], 34, 34, comp1158minVal, comp1158minI, comp1158minJ);
    wire [11:0] comp1159minVal;
    wire [5:0] comp1159minI, comp1159minJ;
    Comparator comp1159(SADValues[2147*12 +: 12], 33, 35, SADValues[2084*12 +: 12], 32, 36, comp1159minVal, comp1159minI, comp1159minJ);
    wire [11:0] comp1160minVal;
    wire [5:0] comp1160minI, comp1160minJ;
    Comparator comp1160(SADValues[2021*12 +: 12], 31, 37, SADValues[1958*12 +: 12], 30, 38, comp1160minVal, comp1160minI, comp1160minJ);
    wire [11:0] comp1161minVal;
    wire [5:0] comp1161minI, comp1161minJ;
    Comparator comp1161(SADValues[1895*12 +: 12], 29, 39, SADValues[1832*12 +: 12], 28, 40, comp1161minVal, comp1161minI, comp1161minJ);
    wire [11:0] comp1162minVal;
    wire [5:0] comp1162minI, comp1162minJ;
    Comparator comp1162(SADValues[1769*12 +: 12], 27, 41, SADValues[1706*12 +: 12], 26, 42, comp1162minVal, comp1162minI, comp1162minJ);
    wire [11:0] comp1163minVal;
    wire [5:0] comp1163minI, comp1163minJ;
    Comparator comp1163(SADValues[1643*12 +: 12], 25, 43, SADValues[1580*12 +: 12], 24, 44, comp1163minVal, comp1163minI, comp1163minJ);
    wire [11:0] comp1164minVal;
    wire [5:0] comp1164minI, comp1164minJ;
    Comparator comp1164(SADValues[1517*12 +: 12], 23, 45, SADValues[1454*12 +: 12], 22, 46, comp1164minVal, comp1164minI, comp1164minJ);
    wire [11:0] comp1165minVal;
    wire [5:0] comp1165minI, comp1165minJ;
    Comparator comp1165(SADValues[1391*12 +: 12], 21, 47, SADValues[1328*12 +: 12], 20, 48, comp1165minVal, comp1165minI, comp1165minJ);
    wire [11:0] comp1166minVal;
    wire [5:0] comp1166minI, comp1166minJ;
    Comparator comp1166(SADValues[1265*12 +: 12], 19, 49, SADValues[1202*12 +: 12], 18, 50, comp1166minVal, comp1166minI, comp1166minJ);
    wire [11:0] comp1167minVal;
    wire [5:0] comp1167minI, comp1167minJ;
    Comparator comp1167(SADValues[1139*12 +: 12], 17, 51, SADValues[1076*12 +: 12], 16, 52, comp1167minVal, comp1167minI, comp1167minJ);
    wire [11:0] comp1168minVal;
    wire [5:0] comp1168minI, comp1168minJ;
    Comparator comp1168(SADValues[1013*12 +: 12], 15, 53, SADValues[950*12 +: 12], 14, 54, comp1168minVal, comp1168minI, comp1168minJ);
    wire [11:0] comp1169minVal;
    wire [5:0] comp1169minI, comp1169minJ;
    Comparator comp1169(SADValues[887*12 +: 12], 13, 55, SADValues[824*12 +: 12], 12, 56, comp1169minVal, comp1169minI, comp1169minJ);
    wire [11:0] comp1170minVal;
    wire [5:0] comp1170minI, comp1170minJ;
    Comparator comp1170(SADValues[761*12 +: 12], 11, 57, SADValues[698*12 +: 12], 10, 58, comp1170minVal, comp1170minI, comp1170minJ);
    wire [11:0] comp1171minVal;
    wire [5:0] comp1171minI, comp1171minJ;
    Comparator comp1171(SADValues[635*12 +: 12], 9, 59, SADValues[572*12 +: 12], 8, 60, comp1171minVal, comp1171minI, comp1171minJ);
    wire [11:0] comp1172minVal;
    wire [5:0] comp1172minI, comp1172minJ;
    Comparator comp1172(SADValues[636*12 +: 12], 9, 60, SADValues[699*12 +: 12], 10, 59, comp1172minVal, comp1172minI, comp1172minJ);
    wire [11:0] comp1173minVal;
    wire [5:0] comp1173minI, comp1173minJ;
    Comparator comp1173(SADValues[762*12 +: 12], 11, 58, SADValues[825*12 +: 12], 12, 57, comp1173minVal, comp1173minI, comp1173minJ);
    wire [11:0] comp1174minVal;
    wire [5:0] comp1174minI, comp1174minJ;
    Comparator comp1174(SADValues[888*12 +: 12], 13, 56, SADValues[951*12 +: 12], 14, 55, comp1174minVal, comp1174minI, comp1174minJ);
    wire [11:0] comp1175minVal;
    wire [5:0] comp1175minI, comp1175minJ;
    Comparator comp1175(SADValues[1014*12 +: 12], 15, 54, SADValues[1077*12 +: 12], 16, 53, comp1175minVal, comp1175minI, comp1175minJ);
    wire [11:0] comp1176minVal;
    wire [5:0] comp1176minI, comp1176minJ;
    Comparator comp1176(SADValues[1140*12 +: 12], 17, 52, SADValues[1203*12 +: 12], 18, 51, comp1176minVal, comp1176minI, comp1176minJ);
    wire [11:0] comp1177minVal;
    wire [5:0] comp1177minI, comp1177minJ;
    Comparator comp1177(SADValues[1266*12 +: 12], 19, 50, SADValues[1329*12 +: 12], 20, 49, comp1177minVal, comp1177minI, comp1177minJ);
    wire [11:0] comp1178minVal;
    wire [5:0] comp1178minI, comp1178minJ;
    Comparator comp1178(SADValues[1392*12 +: 12], 21, 48, SADValues[1455*12 +: 12], 22, 47, comp1178minVal, comp1178minI, comp1178minJ);
    wire [11:0] comp1179minVal;
    wire [5:0] comp1179minI, comp1179minJ;
    Comparator comp1179(SADValues[1518*12 +: 12], 23, 46, SADValues[1581*12 +: 12], 24, 45, comp1179minVal, comp1179minI, comp1179minJ);
    wire [11:0] comp1180minVal;
    wire [5:0] comp1180minI, comp1180minJ;
    Comparator comp1180(SADValues[1644*12 +: 12], 25, 44, SADValues[1707*12 +: 12], 26, 43, comp1180minVal, comp1180minI, comp1180minJ);
    wire [11:0] comp1181minVal;
    wire [5:0] comp1181minI, comp1181minJ;
    Comparator comp1181(SADValues[1770*12 +: 12], 27, 42, SADValues[1833*12 +: 12], 28, 41, comp1181minVal, comp1181minI, comp1181minJ);
    wire [11:0] comp1182minVal;
    wire [5:0] comp1182minI, comp1182minJ;
    Comparator comp1182(SADValues[1896*12 +: 12], 29, 40, SADValues[1959*12 +: 12], 30, 39, comp1182minVal, comp1182minI, comp1182minJ);
    wire [11:0] comp1183minVal;
    wire [5:0] comp1183minI, comp1183minJ;
    Comparator comp1183(SADValues[2022*12 +: 12], 31, 38, SADValues[2085*12 +: 12], 32, 37, comp1183minVal, comp1183minI, comp1183minJ);
    wire [11:0] comp1184minVal;
    wire [5:0] comp1184minI, comp1184minJ;
    Comparator comp1184(SADValues[2148*12 +: 12], 33, 36, SADValues[2211*12 +: 12], 34, 35, comp1184minVal, comp1184minI, comp1184minJ);
    wire [11:0] comp1185minVal;
    wire [5:0] comp1185minI, comp1185minJ;
    Comparator comp1185(SADValues[2274*12 +: 12], 35, 34, SADValues[2337*12 +: 12], 36, 33, comp1185minVal, comp1185minI, comp1185minJ);
    wire [11:0] comp1186minVal;
    wire [5:0] comp1186minI, comp1186minJ;
    Comparator comp1186(SADValues[2400*12 +: 12], 37, 32, SADValues[2463*12 +: 12], 38, 31, comp1186minVal, comp1186minI, comp1186minJ);
    wire [11:0] comp1187minVal;
    wire [5:0] comp1187minI, comp1187minJ;
    Comparator comp1187(SADValues[2526*12 +: 12], 39, 30, SADValues[2589*12 +: 12], 40, 29, comp1187minVal, comp1187minI, comp1187minJ);
    wire [11:0] comp1188minVal;
    wire [5:0] comp1188minI, comp1188minJ;
    Comparator comp1188(SADValues[2652*12 +: 12], 41, 28, SADValues[2715*12 +: 12], 42, 27, comp1188minVal, comp1188minI, comp1188minJ);
    wire [11:0] comp1189minVal;
    wire [5:0] comp1189minI, comp1189minJ;
    Comparator comp1189(SADValues[2778*12 +: 12], 43, 26, SADValues[2841*12 +: 12], 44, 25, comp1189minVal, comp1189minI, comp1189minJ);
    wire [11:0] comp1190minVal;
    wire [5:0] comp1190minI, comp1190minJ;
    Comparator comp1190(SADValues[2904*12 +: 12], 45, 24, SADValues[2967*12 +: 12], 46, 23, comp1190minVal, comp1190minI, comp1190minJ);
    wire [11:0] comp1191minVal;
    wire [5:0] comp1191minI, comp1191minJ;
    Comparator comp1191(SADValues[3030*12 +: 12], 47, 22, SADValues[3093*12 +: 12], 48, 21, comp1191minVal, comp1191minI, comp1191minJ);
    wire [11:0] comp1192minVal;
    wire [5:0] comp1192minI, comp1192minJ;
    Comparator comp1192(SADValues[3156*12 +: 12], 49, 20, SADValues[3219*12 +: 12], 50, 19, comp1192minVal, comp1192minI, comp1192minJ);
    wire [11:0] comp1193minVal;
    wire [5:0] comp1193minI, comp1193minJ;
    Comparator comp1193(SADValues[3282*12 +: 12], 51, 18, SADValues[3345*12 +: 12], 52, 17, comp1193minVal, comp1193minI, comp1193minJ);
    wire [11:0] comp1194minVal;
    wire [5:0] comp1194minI, comp1194minJ;
    Comparator comp1194(SADValues[3408*12 +: 12], 53, 16, SADValues[3471*12 +: 12], 54, 15, comp1194minVal, comp1194minI, comp1194minJ);
    wire [11:0] comp1195minVal;
    wire [5:0] comp1195minI, comp1195minJ;
    Comparator comp1195(SADValues[3534*12 +: 12], 55, 14, SADValues[3597*12 +: 12], 56, 13, comp1195minVal, comp1195minI, comp1195minJ);
    wire [11:0] comp1196minVal;
    wire [5:0] comp1196minI, comp1196minJ;
    Comparator comp1196(SADValues[3660*12 +: 12], 57, 12, SADValues[3723*12 +: 12], 58, 11, comp1196minVal, comp1196minI, comp1196minJ);
    wire [11:0] comp1197minVal;
    wire [5:0] comp1197minI, comp1197minJ;
    Comparator comp1197(SADValues[3786*12 +: 12], 59, 10, SADValues[3849*12 +: 12], 60, 9, comp1197minVal, comp1197minI, comp1197minJ);
    wire [11:0] comp1198minVal;
    wire [5:0] comp1198minI, comp1198minJ;
    Comparator comp1198(SADValues[3850*12 +: 12], 60, 10, SADValues[3787*12 +: 12], 59, 11, comp1198minVal, comp1198minI, comp1198minJ);
    wire [11:0] comp1199minVal;
    wire [5:0] comp1199minI, comp1199minJ;
    Comparator comp1199(SADValues[3724*12 +: 12], 58, 12, SADValues[3661*12 +: 12], 57, 13, comp1199minVal, comp1199minI, comp1199minJ);
    wire [11:0] comp1200minVal;
    wire [5:0] comp1200minI, comp1200minJ;
    Comparator comp1200(SADValues[3598*12 +: 12], 56, 14, SADValues[3535*12 +: 12], 55, 15, comp1200minVal, comp1200minI, comp1200minJ);
    wire [11:0] comp1201minVal;
    wire [5:0] comp1201minI, comp1201minJ;
    Comparator comp1201(SADValues[3472*12 +: 12], 54, 16, SADValues[3409*12 +: 12], 53, 17, comp1201minVal, comp1201minI, comp1201minJ);
    wire [11:0] comp1202minVal;
    wire [5:0] comp1202minI, comp1202minJ;
    Comparator comp1202(SADValues[3346*12 +: 12], 52, 18, SADValues[3283*12 +: 12], 51, 19, comp1202minVal, comp1202minI, comp1202minJ);
    wire [11:0] comp1203minVal;
    wire [5:0] comp1203minI, comp1203minJ;
    Comparator comp1203(SADValues[3220*12 +: 12], 50, 20, SADValues[3157*12 +: 12], 49, 21, comp1203minVal, comp1203minI, comp1203minJ);
    wire [11:0] comp1204minVal;
    wire [5:0] comp1204minI, comp1204minJ;
    Comparator comp1204(SADValues[3094*12 +: 12], 48, 22, SADValues[3031*12 +: 12], 47, 23, comp1204minVal, comp1204minI, comp1204minJ);
    wire [11:0] comp1205minVal;
    wire [5:0] comp1205minI, comp1205minJ;
    Comparator comp1205(SADValues[2968*12 +: 12], 46, 24, SADValues[2905*12 +: 12], 45, 25, comp1205minVal, comp1205minI, comp1205minJ);
    wire [11:0] comp1206minVal;
    wire [5:0] comp1206minI, comp1206minJ;
    Comparator comp1206(SADValues[2842*12 +: 12], 44, 26, SADValues[2779*12 +: 12], 43, 27, comp1206minVal, comp1206minI, comp1206minJ);
    wire [11:0] comp1207minVal;
    wire [5:0] comp1207minI, comp1207minJ;
    Comparator comp1207(SADValues[2716*12 +: 12], 42, 28, SADValues[2653*12 +: 12], 41, 29, comp1207minVal, comp1207minI, comp1207minJ);
    wire [11:0] comp1208minVal;
    wire [5:0] comp1208minI, comp1208minJ;
    Comparator comp1208(SADValues[2590*12 +: 12], 40, 30, SADValues[2527*12 +: 12], 39, 31, comp1208minVal, comp1208minI, comp1208minJ);
    wire [11:0] comp1209minVal;
    wire [5:0] comp1209minI, comp1209minJ;
    Comparator comp1209(SADValues[2464*12 +: 12], 38, 32, SADValues[2401*12 +: 12], 37, 33, comp1209minVal, comp1209minI, comp1209minJ);
    wire [11:0] comp1210minVal;
    wire [5:0] comp1210minI, comp1210minJ;
    Comparator comp1210(SADValues[2338*12 +: 12], 36, 34, SADValues[2275*12 +: 12], 35, 35, comp1210minVal, comp1210minI, comp1210minJ);
    wire [11:0] comp1211minVal;
    wire [5:0] comp1211minI, comp1211minJ;
    Comparator comp1211(SADValues[2212*12 +: 12], 34, 36, SADValues[2149*12 +: 12], 33, 37, comp1211minVal, comp1211minI, comp1211minJ);
    wire [11:0] comp1212minVal;
    wire [5:0] comp1212minI, comp1212minJ;
    Comparator comp1212(SADValues[2086*12 +: 12], 32, 38, SADValues[2023*12 +: 12], 31, 39, comp1212minVal, comp1212minI, comp1212minJ);
    wire [11:0] comp1213minVal;
    wire [5:0] comp1213minI, comp1213minJ;
    Comparator comp1213(SADValues[1960*12 +: 12], 30, 40, SADValues[1897*12 +: 12], 29, 41, comp1213minVal, comp1213minI, comp1213minJ);
    wire [11:0] comp1214minVal;
    wire [5:0] comp1214minI, comp1214minJ;
    Comparator comp1214(SADValues[1834*12 +: 12], 28, 42, SADValues[1771*12 +: 12], 27, 43, comp1214minVal, comp1214minI, comp1214minJ);
    wire [11:0] comp1215minVal;
    wire [5:0] comp1215minI, comp1215minJ;
    Comparator comp1215(SADValues[1708*12 +: 12], 26, 44, SADValues[1645*12 +: 12], 25, 45, comp1215minVal, comp1215minI, comp1215minJ);
    wire [11:0] comp1216minVal;
    wire [5:0] comp1216minI, comp1216minJ;
    Comparator comp1216(SADValues[1582*12 +: 12], 24, 46, SADValues[1519*12 +: 12], 23, 47, comp1216minVal, comp1216minI, comp1216minJ);
    wire [11:0] comp1217minVal;
    wire [5:0] comp1217minI, comp1217minJ;
    Comparator comp1217(SADValues[1456*12 +: 12], 22, 48, SADValues[1393*12 +: 12], 21, 49, comp1217minVal, comp1217minI, comp1217minJ);
    wire [11:0] comp1218minVal;
    wire [5:0] comp1218minI, comp1218minJ;
    Comparator comp1218(SADValues[1330*12 +: 12], 20, 50, SADValues[1267*12 +: 12], 19, 51, comp1218minVal, comp1218minI, comp1218minJ);
    wire [11:0] comp1219minVal;
    wire [5:0] comp1219minI, comp1219minJ;
    Comparator comp1219(SADValues[1204*12 +: 12], 18, 52, SADValues[1141*12 +: 12], 17, 53, comp1219minVal, comp1219minI, comp1219minJ);
    wire [11:0] comp1220minVal;
    wire [5:0] comp1220minI, comp1220minJ;
    Comparator comp1220(SADValues[1078*12 +: 12], 16, 54, SADValues[1015*12 +: 12], 15, 55, comp1220minVal, comp1220minI, comp1220minJ);
    wire [11:0] comp1221minVal;
    wire [5:0] comp1221minI, comp1221minJ;
    Comparator comp1221(SADValues[952*12 +: 12], 14, 56, SADValues[889*12 +: 12], 13, 57, comp1221minVal, comp1221minI, comp1221minJ);
    wire [11:0] comp1222minVal;
    wire [5:0] comp1222minI, comp1222minJ;
    Comparator comp1222(SADValues[826*12 +: 12], 12, 58, SADValues[763*12 +: 12], 11, 59, comp1222minVal, comp1222minI, comp1222minJ);
    wire [11:0] comp1223minVal;
    wire [5:0] comp1223minI, comp1223minJ;
    Comparator comp1223(SADValues[700*12 +: 12], 10, 60, SADValues[764*12 +: 12], 11, 60, comp1223minVal, comp1223minI, comp1223minJ);
    wire [11:0] comp1224minVal;
    wire [5:0] comp1224minI, comp1224minJ;
    Comparator comp1224(SADValues[827*12 +: 12], 12, 59, SADValues[890*12 +: 12], 13, 58, comp1224minVal, comp1224minI, comp1224minJ);
    wire [11:0] comp1225minVal;
    wire [5:0] comp1225minI, comp1225minJ;
    Comparator comp1225(SADValues[953*12 +: 12], 14, 57, SADValues[1016*12 +: 12], 15, 56, comp1225minVal, comp1225minI, comp1225minJ);
    wire [11:0] comp1226minVal;
    wire [5:0] comp1226minI, comp1226minJ;
    Comparator comp1226(SADValues[1079*12 +: 12], 16, 55, SADValues[1142*12 +: 12], 17, 54, comp1226minVal, comp1226minI, comp1226minJ);
    wire [11:0] comp1227minVal;
    wire [5:0] comp1227minI, comp1227minJ;
    Comparator comp1227(SADValues[1205*12 +: 12], 18, 53, SADValues[1268*12 +: 12], 19, 52, comp1227minVal, comp1227minI, comp1227minJ);
    wire [11:0] comp1228minVal;
    wire [5:0] comp1228minI, comp1228minJ;
    Comparator comp1228(SADValues[1331*12 +: 12], 20, 51, SADValues[1394*12 +: 12], 21, 50, comp1228minVal, comp1228minI, comp1228minJ);
    wire [11:0] comp1229minVal;
    wire [5:0] comp1229minI, comp1229minJ;
    Comparator comp1229(SADValues[1457*12 +: 12], 22, 49, SADValues[1520*12 +: 12], 23, 48, comp1229minVal, comp1229minI, comp1229minJ);
    wire [11:0] comp1230minVal;
    wire [5:0] comp1230minI, comp1230minJ;
    Comparator comp1230(SADValues[1583*12 +: 12], 24, 47, SADValues[1646*12 +: 12], 25, 46, comp1230minVal, comp1230minI, comp1230minJ);
    wire [11:0] comp1231minVal;
    wire [5:0] comp1231minI, comp1231minJ;
    Comparator comp1231(SADValues[1709*12 +: 12], 26, 45, SADValues[1772*12 +: 12], 27, 44, comp1231minVal, comp1231minI, comp1231minJ);
    wire [11:0] comp1232minVal;
    wire [5:0] comp1232minI, comp1232minJ;
    Comparator comp1232(SADValues[1835*12 +: 12], 28, 43, SADValues[1898*12 +: 12], 29, 42, comp1232minVal, comp1232minI, comp1232minJ);
    wire [11:0] comp1233minVal;
    wire [5:0] comp1233minI, comp1233minJ;
    Comparator comp1233(SADValues[1961*12 +: 12], 30, 41, SADValues[2024*12 +: 12], 31, 40, comp1233minVal, comp1233minI, comp1233minJ);
    wire [11:0] comp1234minVal;
    wire [5:0] comp1234minI, comp1234minJ;
    Comparator comp1234(SADValues[2087*12 +: 12], 32, 39, SADValues[2150*12 +: 12], 33, 38, comp1234minVal, comp1234minI, comp1234minJ);
    wire [11:0] comp1235minVal;
    wire [5:0] comp1235minI, comp1235minJ;
    Comparator comp1235(SADValues[2213*12 +: 12], 34, 37, SADValues[2276*12 +: 12], 35, 36, comp1235minVal, comp1235minI, comp1235minJ);
    wire [11:0] comp1236minVal;
    wire [5:0] comp1236minI, comp1236minJ;
    Comparator comp1236(SADValues[2339*12 +: 12], 36, 35, SADValues[2402*12 +: 12], 37, 34, comp1236minVal, comp1236minI, comp1236minJ);
    wire [11:0] comp1237minVal;
    wire [5:0] comp1237minI, comp1237minJ;
    Comparator comp1237(SADValues[2465*12 +: 12], 38, 33, SADValues[2528*12 +: 12], 39, 32, comp1237minVal, comp1237minI, comp1237minJ);
    wire [11:0] comp1238minVal;
    wire [5:0] comp1238minI, comp1238minJ;
    Comparator comp1238(SADValues[2591*12 +: 12], 40, 31, SADValues[2654*12 +: 12], 41, 30, comp1238minVal, comp1238minI, comp1238minJ);
    wire [11:0] comp1239minVal;
    wire [5:0] comp1239minI, comp1239minJ;
    Comparator comp1239(SADValues[2717*12 +: 12], 42, 29, SADValues[2780*12 +: 12], 43, 28, comp1239minVal, comp1239minI, comp1239minJ);
    wire [11:0] comp1240minVal;
    wire [5:0] comp1240minI, comp1240minJ;
    Comparator comp1240(SADValues[2843*12 +: 12], 44, 27, SADValues[2906*12 +: 12], 45, 26, comp1240minVal, comp1240minI, comp1240minJ);
    wire [11:0] comp1241minVal;
    wire [5:0] comp1241minI, comp1241minJ;
    Comparator comp1241(SADValues[2969*12 +: 12], 46, 25, SADValues[3032*12 +: 12], 47, 24, comp1241minVal, comp1241minI, comp1241minJ);
    wire [11:0] comp1242minVal;
    wire [5:0] comp1242minI, comp1242minJ;
    Comparator comp1242(SADValues[3095*12 +: 12], 48, 23, SADValues[3158*12 +: 12], 49, 22, comp1242minVal, comp1242minI, comp1242minJ);
    wire [11:0] comp1243minVal;
    wire [5:0] comp1243minI, comp1243minJ;
    Comparator comp1243(SADValues[3221*12 +: 12], 50, 21, SADValues[3284*12 +: 12], 51, 20, comp1243minVal, comp1243minI, comp1243minJ);
    wire [11:0] comp1244minVal;
    wire [5:0] comp1244minI, comp1244minJ;
    Comparator comp1244(SADValues[3347*12 +: 12], 52, 19, SADValues[3410*12 +: 12], 53, 18, comp1244minVal, comp1244minI, comp1244minJ);
    wire [11:0] comp1245minVal;
    wire [5:0] comp1245minI, comp1245minJ;
    Comparator comp1245(SADValues[3473*12 +: 12], 54, 17, SADValues[3536*12 +: 12], 55, 16, comp1245minVal, comp1245minI, comp1245minJ);
    wire [11:0] comp1246minVal;
    wire [5:0] comp1246minI, comp1246minJ;
    Comparator comp1246(SADValues[3599*12 +: 12], 56, 15, SADValues[3662*12 +: 12], 57, 14, comp1246minVal, comp1246minI, comp1246minJ);
    wire [11:0] comp1247minVal;
    wire [5:0] comp1247minI, comp1247minJ;
    Comparator comp1247(SADValues[3725*12 +: 12], 58, 13, SADValues[3788*12 +: 12], 59, 12, comp1247minVal, comp1247minI, comp1247minJ);
    wire [11:0] comp1248minVal;
    wire [5:0] comp1248minI, comp1248minJ;
    Comparator comp1248(SADValues[3851*12 +: 12], 60, 11, SADValues[3852*12 +: 12], 60, 12, comp1248minVal, comp1248minI, comp1248minJ);
    wire [11:0] comp1249minVal;
    wire [5:0] comp1249minI, comp1249minJ;
    Comparator comp1249(SADValues[3789*12 +: 12], 59, 13, SADValues[3726*12 +: 12], 58, 14, comp1249minVal, comp1249minI, comp1249minJ);
    wire [11:0] comp1250minVal;
    wire [5:0] comp1250minI, comp1250minJ;
    Comparator comp1250(SADValues[3663*12 +: 12], 57, 15, SADValues[3600*12 +: 12], 56, 16, comp1250minVal, comp1250minI, comp1250minJ);
    wire [11:0] comp1251minVal;
    wire [5:0] comp1251minI, comp1251minJ;
    Comparator comp1251(SADValues[3537*12 +: 12], 55, 17, SADValues[3474*12 +: 12], 54, 18, comp1251minVal, comp1251minI, comp1251minJ);
    wire [11:0] comp1252minVal;
    wire [5:0] comp1252minI, comp1252minJ;
    Comparator comp1252(SADValues[3411*12 +: 12], 53, 19, SADValues[3348*12 +: 12], 52, 20, comp1252minVal, comp1252minI, comp1252minJ);
    wire [11:0] comp1253minVal;
    wire [5:0] comp1253minI, comp1253minJ;
    Comparator comp1253(SADValues[3285*12 +: 12], 51, 21, SADValues[3222*12 +: 12], 50, 22, comp1253minVal, comp1253minI, comp1253minJ);
    wire [11:0] comp1254minVal;
    wire [5:0] comp1254minI, comp1254minJ;
    Comparator comp1254(SADValues[3159*12 +: 12], 49, 23, SADValues[3096*12 +: 12], 48, 24, comp1254minVal, comp1254minI, comp1254minJ);
    wire [11:0] comp1255minVal;
    wire [5:0] comp1255minI, comp1255minJ;
    Comparator comp1255(SADValues[3033*12 +: 12], 47, 25, SADValues[2970*12 +: 12], 46, 26, comp1255minVal, comp1255minI, comp1255minJ);
    wire [11:0] comp1256minVal;
    wire [5:0] comp1256minI, comp1256minJ;
    Comparator comp1256(SADValues[2907*12 +: 12], 45, 27, SADValues[2844*12 +: 12], 44, 28, comp1256minVal, comp1256minI, comp1256minJ);
    wire [11:0] comp1257minVal;
    wire [5:0] comp1257minI, comp1257minJ;
    Comparator comp1257(SADValues[2781*12 +: 12], 43, 29, SADValues[2718*12 +: 12], 42, 30, comp1257minVal, comp1257minI, comp1257minJ);
    wire [11:0] comp1258minVal;
    wire [5:0] comp1258minI, comp1258minJ;
    Comparator comp1258(SADValues[2655*12 +: 12], 41, 31, SADValues[2592*12 +: 12], 40, 32, comp1258minVal, comp1258minI, comp1258minJ);
    wire [11:0] comp1259minVal;
    wire [5:0] comp1259minI, comp1259minJ;
    Comparator comp1259(SADValues[2529*12 +: 12], 39, 33, SADValues[2466*12 +: 12], 38, 34, comp1259minVal, comp1259minI, comp1259minJ);
    wire [11:0] comp1260minVal;
    wire [5:0] comp1260minI, comp1260minJ;
    Comparator comp1260(SADValues[2403*12 +: 12], 37, 35, SADValues[2340*12 +: 12], 36, 36, comp1260minVal, comp1260minI, comp1260minJ);
    wire [11:0] comp1261minVal;
    wire [5:0] comp1261minI, comp1261minJ;
    Comparator comp1261(SADValues[2277*12 +: 12], 35, 37, SADValues[2214*12 +: 12], 34, 38, comp1261minVal, comp1261minI, comp1261minJ);
    wire [11:0] comp1262minVal;
    wire [5:0] comp1262minI, comp1262minJ;
    Comparator comp1262(SADValues[2151*12 +: 12], 33, 39, SADValues[2088*12 +: 12], 32, 40, comp1262minVal, comp1262minI, comp1262minJ);
    wire [11:0] comp1263minVal;
    wire [5:0] comp1263minI, comp1263minJ;
    Comparator comp1263(SADValues[2025*12 +: 12], 31, 41, SADValues[1962*12 +: 12], 30, 42, comp1263minVal, comp1263minI, comp1263minJ);
    wire [11:0] comp1264minVal;
    wire [5:0] comp1264minI, comp1264minJ;
    Comparator comp1264(SADValues[1899*12 +: 12], 29, 43, SADValues[1836*12 +: 12], 28, 44, comp1264minVal, comp1264minI, comp1264minJ);
    wire [11:0] comp1265minVal;
    wire [5:0] comp1265minI, comp1265minJ;
    Comparator comp1265(SADValues[1773*12 +: 12], 27, 45, SADValues[1710*12 +: 12], 26, 46, comp1265minVal, comp1265minI, comp1265minJ);
    wire [11:0] comp1266minVal;
    wire [5:0] comp1266minI, comp1266minJ;
    Comparator comp1266(SADValues[1647*12 +: 12], 25, 47, SADValues[1584*12 +: 12], 24, 48, comp1266minVal, comp1266minI, comp1266minJ);
    wire [11:0] comp1267minVal;
    wire [5:0] comp1267minI, comp1267minJ;
    Comparator comp1267(SADValues[1521*12 +: 12], 23, 49, SADValues[1458*12 +: 12], 22, 50, comp1267minVal, comp1267minI, comp1267minJ);
    wire [11:0] comp1268minVal;
    wire [5:0] comp1268minI, comp1268minJ;
    Comparator comp1268(SADValues[1395*12 +: 12], 21, 51, SADValues[1332*12 +: 12], 20, 52, comp1268minVal, comp1268minI, comp1268minJ);
    wire [11:0] comp1269minVal;
    wire [5:0] comp1269minI, comp1269minJ;
    Comparator comp1269(SADValues[1269*12 +: 12], 19, 53, SADValues[1206*12 +: 12], 18, 54, comp1269minVal, comp1269minI, comp1269minJ);
    wire [11:0] comp1270minVal;
    wire [5:0] comp1270minI, comp1270minJ;
    Comparator comp1270(SADValues[1143*12 +: 12], 17, 55, SADValues[1080*12 +: 12], 16, 56, comp1270minVal, comp1270minI, comp1270minJ);
    wire [11:0] comp1271minVal;
    wire [5:0] comp1271minI, comp1271minJ;
    Comparator comp1271(SADValues[1017*12 +: 12], 15, 57, SADValues[954*12 +: 12], 14, 58, comp1271minVal, comp1271minI, comp1271minJ);
    wire [11:0] comp1272minVal;
    wire [5:0] comp1272minI, comp1272minJ;
    Comparator comp1272(SADValues[891*12 +: 12], 13, 59, SADValues[828*12 +: 12], 12, 60, comp1272minVal, comp1272minI, comp1272minJ);
    wire [11:0] comp1273minVal;
    wire [5:0] comp1273minI, comp1273minJ;
    Comparator comp1273(SADValues[892*12 +: 12], 13, 60, SADValues[955*12 +: 12], 14, 59, comp1273minVal, comp1273minI, comp1273minJ);
    wire [11:0] comp1274minVal;
    wire [5:0] comp1274minI, comp1274minJ;
    Comparator comp1274(SADValues[1018*12 +: 12], 15, 58, SADValues[1081*12 +: 12], 16, 57, comp1274minVal, comp1274minI, comp1274minJ);
    wire [11:0] comp1275minVal;
    wire [5:0] comp1275minI, comp1275minJ;
    Comparator comp1275(SADValues[1144*12 +: 12], 17, 56, SADValues[1207*12 +: 12], 18, 55, comp1275minVal, comp1275minI, comp1275minJ);
    wire [11:0] comp1276minVal;
    wire [5:0] comp1276minI, comp1276minJ;
    Comparator comp1276(SADValues[1270*12 +: 12], 19, 54, SADValues[1333*12 +: 12], 20, 53, comp1276minVal, comp1276minI, comp1276minJ);
    wire [11:0] comp1277minVal;
    wire [5:0] comp1277minI, comp1277minJ;
    Comparator comp1277(SADValues[1396*12 +: 12], 21, 52, SADValues[1459*12 +: 12], 22, 51, comp1277minVal, comp1277minI, comp1277minJ);
    wire [11:0] comp1278minVal;
    wire [5:0] comp1278minI, comp1278minJ;
    Comparator comp1278(SADValues[1522*12 +: 12], 23, 50, SADValues[1585*12 +: 12], 24, 49, comp1278minVal, comp1278minI, comp1278minJ);
    wire [11:0] comp1279minVal;
    wire [5:0] comp1279minI, comp1279minJ;
    Comparator comp1279(SADValues[1648*12 +: 12], 25, 48, SADValues[1711*12 +: 12], 26, 47, comp1279minVal, comp1279minI, comp1279minJ);
    wire [11:0] comp1280minVal;
    wire [5:0] comp1280minI, comp1280minJ;
    Comparator comp1280(SADValues[1774*12 +: 12], 27, 46, SADValues[1837*12 +: 12], 28, 45, comp1280minVal, comp1280minI, comp1280minJ);
    wire [11:0] comp1281minVal;
    wire [5:0] comp1281minI, comp1281minJ;
    Comparator comp1281(SADValues[1900*12 +: 12], 29, 44, SADValues[1963*12 +: 12], 30, 43, comp1281minVal, comp1281minI, comp1281minJ);
    wire [11:0] comp1282minVal;
    wire [5:0] comp1282minI, comp1282minJ;
    Comparator comp1282(SADValues[2026*12 +: 12], 31, 42, SADValues[2089*12 +: 12], 32, 41, comp1282minVal, comp1282minI, comp1282minJ);
    wire [11:0] comp1283minVal;
    wire [5:0] comp1283minI, comp1283minJ;
    Comparator comp1283(SADValues[2152*12 +: 12], 33, 40, SADValues[2215*12 +: 12], 34, 39, comp1283minVal, comp1283minI, comp1283minJ);
    wire [11:0] comp1284minVal;
    wire [5:0] comp1284minI, comp1284minJ;
    Comparator comp1284(SADValues[2278*12 +: 12], 35, 38, SADValues[2341*12 +: 12], 36, 37, comp1284minVal, comp1284minI, comp1284minJ);
    wire [11:0] comp1285minVal;
    wire [5:0] comp1285minI, comp1285minJ;
    Comparator comp1285(SADValues[2404*12 +: 12], 37, 36, SADValues[2467*12 +: 12], 38, 35, comp1285minVal, comp1285minI, comp1285minJ);
    wire [11:0] comp1286minVal;
    wire [5:0] comp1286minI, comp1286minJ;
    Comparator comp1286(SADValues[2530*12 +: 12], 39, 34, SADValues[2593*12 +: 12], 40, 33, comp1286minVal, comp1286minI, comp1286minJ);
    wire [11:0] comp1287minVal;
    wire [5:0] comp1287minI, comp1287minJ;
    Comparator comp1287(SADValues[2656*12 +: 12], 41, 32, SADValues[2719*12 +: 12], 42, 31, comp1287minVal, comp1287minI, comp1287minJ);
    wire [11:0] comp1288minVal;
    wire [5:0] comp1288minI, comp1288minJ;
    Comparator comp1288(SADValues[2782*12 +: 12], 43, 30, SADValues[2845*12 +: 12], 44, 29, comp1288minVal, comp1288minI, comp1288minJ);
    wire [11:0] comp1289minVal;
    wire [5:0] comp1289minI, comp1289minJ;
    Comparator comp1289(SADValues[2908*12 +: 12], 45, 28, SADValues[2971*12 +: 12], 46, 27, comp1289minVal, comp1289minI, comp1289minJ);
    wire [11:0] comp1290minVal;
    wire [5:0] comp1290minI, comp1290minJ;
    Comparator comp1290(SADValues[3034*12 +: 12], 47, 26, SADValues[3097*12 +: 12], 48, 25, comp1290minVal, comp1290minI, comp1290minJ);
    wire [11:0] comp1291minVal;
    wire [5:0] comp1291minI, comp1291minJ;
    Comparator comp1291(SADValues[3160*12 +: 12], 49, 24, SADValues[3223*12 +: 12], 50, 23, comp1291minVal, comp1291minI, comp1291minJ);
    wire [11:0] comp1292minVal;
    wire [5:0] comp1292minI, comp1292minJ;
    Comparator comp1292(SADValues[3286*12 +: 12], 51, 22, SADValues[3349*12 +: 12], 52, 21, comp1292minVal, comp1292minI, comp1292minJ);
    wire [11:0] comp1293minVal;
    wire [5:0] comp1293minI, comp1293minJ;
    Comparator comp1293(SADValues[3412*12 +: 12], 53, 20, SADValues[3475*12 +: 12], 54, 19, comp1293minVal, comp1293minI, comp1293minJ);
    wire [11:0] comp1294minVal;
    wire [5:0] comp1294minI, comp1294minJ;
    Comparator comp1294(SADValues[3538*12 +: 12], 55, 18, SADValues[3601*12 +: 12], 56, 17, comp1294minVal, comp1294minI, comp1294minJ);
    wire [11:0] comp1295minVal;
    wire [5:0] comp1295minI, comp1295minJ;
    Comparator comp1295(SADValues[3664*12 +: 12], 57, 16, SADValues[3727*12 +: 12], 58, 15, comp1295minVal, comp1295minI, comp1295minJ);
    wire [11:0] comp1296minVal;
    wire [5:0] comp1296minI, comp1296minJ;
    Comparator comp1296(SADValues[3790*12 +: 12], 59, 14, SADValues[3853*12 +: 12], 60, 13, comp1296minVal, comp1296minI, comp1296minJ);
    wire [11:0] comp1297minVal;
    wire [5:0] comp1297minI, comp1297minJ;
    Comparator comp1297(SADValues[3854*12 +: 12], 60, 14, SADValues[3791*12 +: 12], 59, 15, comp1297minVal, comp1297minI, comp1297minJ);
    wire [11:0] comp1298minVal;
    wire [5:0] comp1298minI, comp1298minJ;
    Comparator comp1298(SADValues[3728*12 +: 12], 58, 16, SADValues[3665*12 +: 12], 57, 17, comp1298minVal, comp1298minI, comp1298minJ);
    wire [11:0] comp1299minVal;
    wire [5:0] comp1299minI, comp1299minJ;
    Comparator comp1299(SADValues[3602*12 +: 12], 56, 18, SADValues[3539*12 +: 12], 55, 19, comp1299minVal, comp1299minI, comp1299minJ);
    wire [11:0] comp1300minVal;
    wire [5:0] comp1300minI, comp1300minJ;
    Comparator comp1300(SADValues[3476*12 +: 12], 54, 20, SADValues[3413*12 +: 12], 53, 21, comp1300minVal, comp1300minI, comp1300minJ);
    wire [11:0] comp1301minVal;
    wire [5:0] comp1301minI, comp1301minJ;
    Comparator comp1301(SADValues[3350*12 +: 12], 52, 22, SADValues[3287*12 +: 12], 51, 23, comp1301minVal, comp1301minI, comp1301minJ);
    wire [11:0] comp1302minVal;
    wire [5:0] comp1302minI, comp1302minJ;
    Comparator comp1302(SADValues[3224*12 +: 12], 50, 24, SADValues[3161*12 +: 12], 49, 25, comp1302minVal, comp1302minI, comp1302minJ);
    wire [11:0] comp1303minVal;
    wire [5:0] comp1303minI, comp1303minJ;
    Comparator comp1303(SADValues[3098*12 +: 12], 48, 26, SADValues[3035*12 +: 12], 47, 27, comp1303minVal, comp1303minI, comp1303minJ);
    wire [11:0] comp1304minVal;
    wire [5:0] comp1304minI, comp1304minJ;
    Comparator comp1304(SADValues[2972*12 +: 12], 46, 28, SADValues[2909*12 +: 12], 45, 29, comp1304minVal, comp1304minI, comp1304minJ);
    wire [11:0] comp1305minVal;
    wire [5:0] comp1305minI, comp1305minJ;
    Comparator comp1305(SADValues[2846*12 +: 12], 44, 30, SADValues[2783*12 +: 12], 43, 31, comp1305minVal, comp1305minI, comp1305minJ);
    wire [11:0] comp1306minVal;
    wire [5:0] comp1306minI, comp1306minJ;
    Comparator comp1306(SADValues[2720*12 +: 12], 42, 32, SADValues[2657*12 +: 12], 41, 33, comp1306minVal, comp1306minI, comp1306minJ);
    wire [11:0] comp1307minVal;
    wire [5:0] comp1307minI, comp1307minJ;
    Comparator comp1307(SADValues[2594*12 +: 12], 40, 34, SADValues[2531*12 +: 12], 39, 35, comp1307minVal, comp1307minI, comp1307minJ);
    wire [11:0] comp1308minVal;
    wire [5:0] comp1308minI, comp1308minJ;
    Comparator comp1308(SADValues[2468*12 +: 12], 38, 36, SADValues[2405*12 +: 12], 37, 37, comp1308minVal, comp1308minI, comp1308minJ);
    wire [11:0] comp1309minVal;
    wire [5:0] comp1309minI, comp1309minJ;
    Comparator comp1309(SADValues[2342*12 +: 12], 36, 38, SADValues[2279*12 +: 12], 35, 39, comp1309minVal, comp1309minI, comp1309minJ);
    wire [11:0] comp1310minVal;
    wire [5:0] comp1310minI, comp1310minJ;
    Comparator comp1310(SADValues[2216*12 +: 12], 34, 40, SADValues[2153*12 +: 12], 33, 41, comp1310minVal, comp1310minI, comp1310minJ);
    wire [11:0] comp1311minVal;
    wire [5:0] comp1311minI, comp1311minJ;
    Comparator comp1311(SADValues[2090*12 +: 12], 32, 42, SADValues[2027*12 +: 12], 31, 43, comp1311minVal, comp1311minI, comp1311minJ);
    wire [11:0] comp1312minVal;
    wire [5:0] comp1312minI, comp1312minJ;
    Comparator comp1312(SADValues[1964*12 +: 12], 30, 44, SADValues[1901*12 +: 12], 29, 45, comp1312minVal, comp1312minI, comp1312minJ);
    wire [11:0] comp1313minVal;
    wire [5:0] comp1313minI, comp1313minJ;
    Comparator comp1313(SADValues[1838*12 +: 12], 28, 46, SADValues[1775*12 +: 12], 27, 47, comp1313minVal, comp1313minI, comp1313minJ);
    wire [11:0] comp1314minVal;
    wire [5:0] comp1314minI, comp1314minJ;
    Comparator comp1314(SADValues[1712*12 +: 12], 26, 48, SADValues[1649*12 +: 12], 25, 49, comp1314minVal, comp1314minI, comp1314minJ);
    wire [11:0] comp1315minVal;
    wire [5:0] comp1315minI, comp1315minJ;
    Comparator comp1315(SADValues[1586*12 +: 12], 24, 50, SADValues[1523*12 +: 12], 23, 51, comp1315minVal, comp1315minI, comp1315minJ);
    wire [11:0] comp1316minVal;
    wire [5:0] comp1316minI, comp1316minJ;
    Comparator comp1316(SADValues[1460*12 +: 12], 22, 52, SADValues[1397*12 +: 12], 21, 53, comp1316minVal, comp1316minI, comp1316minJ);
    wire [11:0] comp1317minVal;
    wire [5:0] comp1317minI, comp1317minJ;
    Comparator comp1317(SADValues[1334*12 +: 12], 20, 54, SADValues[1271*12 +: 12], 19, 55, comp1317minVal, comp1317minI, comp1317minJ);
    wire [11:0] comp1318minVal;
    wire [5:0] comp1318minI, comp1318minJ;
    Comparator comp1318(SADValues[1208*12 +: 12], 18, 56, SADValues[1145*12 +: 12], 17, 57, comp1318minVal, comp1318minI, comp1318minJ);
    wire [11:0] comp1319minVal;
    wire [5:0] comp1319minI, comp1319minJ;
    Comparator comp1319(SADValues[1082*12 +: 12], 16, 58, SADValues[1019*12 +: 12], 15, 59, comp1319minVal, comp1319minI, comp1319minJ);
    wire [11:0] comp1320minVal;
    wire [5:0] comp1320minI, comp1320minJ;
    Comparator comp1320(SADValues[956*12 +: 12], 14, 60, SADValues[1020*12 +: 12], 15, 60, comp1320minVal, comp1320minI, comp1320minJ);
    wire [11:0] comp1321minVal;
    wire [5:0] comp1321minI, comp1321minJ;
    Comparator comp1321(SADValues[1083*12 +: 12], 16, 59, SADValues[1146*12 +: 12], 17, 58, comp1321minVal, comp1321minI, comp1321minJ);
    wire [11:0] comp1322minVal;
    wire [5:0] comp1322minI, comp1322minJ;
    Comparator comp1322(SADValues[1209*12 +: 12], 18, 57, SADValues[1272*12 +: 12], 19, 56, comp1322minVal, comp1322minI, comp1322minJ);
    wire [11:0] comp1323minVal;
    wire [5:0] comp1323minI, comp1323minJ;
    Comparator comp1323(SADValues[1335*12 +: 12], 20, 55, SADValues[1398*12 +: 12], 21, 54, comp1323minVal, comp1323minI, comp1323minJ);
    wire [11:0] comp1324minVal;
    wire [5:0] comp1324minI, comp1324minJ;
    Comparator comp1324(SADValues[1461*12 +: 12], 22, 53, SADValues[1524*12 +: 12], 23, 52, comp1324minVal, comp1324minI, comp1324minJ);
    wire [11:0] comp1325minVal;
    wire [5:0] comp1325minI, comp1325minJ;
    Comparator comp1325(SADValues[1587*12 +: 12], 24, 51, SADValues[1650*12 +: 12], 25, 50, comp1325minVal, comp1325minI, comp1325minJ);
    wire [11:0] comp1326minVal;
    wire [5:0] comp1326minI, comp1326minJ;
    Comparator comp1326(SADValues[1713*12 +: 12], 26, 49, SADValues[1776*12 +: 12], 27, 48, comp1326minVal, comp1326minI, comp1326minJ);
    wire [11:0] comp1327minVal;
    wire [5:0] comp1327minI, comp1327minJ;
    Comparator comp1327(SADValues[1839*12 +: 12], 28, 47, SADValues[1902*12 +: 12], 29, 46, comp1327minVal, comp1327minI, comp1327minJ);
    wire [11:0] comp1328minVal;
    wire [5:0] comp1328minI, comp1328minJ;
    Comparator comp1328(SADValues[1965*12 +: 12], 30, 45, SADValues[2028*12 +: 12], 31, 44, comp1328minVal, comp1328minI, comp1328minJ);
    wire [11:0] comp1329minVal;
    wire [5:0] comp1329minI, comp1329minJ;
    Comparator comp1329(SADValues[2091*12 +: 12], 32, 43, SADValues[2154*12 +: 12], 33, 42, comp1329minVal, comp1329minI, comp1329minJ);
    wire [11:0] comp1330minVal;
    wire [5:0] comp1330minI, comp1330minJ;
    Comparator comp1330(SADValues[2217*12 +: 12], 34, 41, SADValues[2280*12 +: 12], 35, 40, comp1330minVal, comp1330minI, comp1330minJ);
    wire [11:0] comp1331minVal;
    wire [5:0] comp1331minI, comp1331minJ;
    Comparator comp1331(SADValues[2343*12 +: 12], 36, 39, SADValues[2406*12 +: 12], 37, 38, comp1331minVal, comp1331minI, comp1331minJ);
    wire [11:0] comp1332minVal;
    wire [5:0] comp1332minI, comp1332minJ;
    Comparator comp1332(SADValues[2469*12 +: 12], 38, 37, SADValues[2532*12 +: 12], 39, 36, comp1332minVal, comp1332minI, comp1332minJ);
    wire [11:0] comp1333minVal;
    wire [5:0] comp1333minI, comp1333minJ;
    Comparator comp1333(SADValues[2595*12 +: 12], 40, 35, SADValues[2658*12 +: 12], 41, 34, comp1333minVal, comp1333minI, comp1333minJ);
    wire [11:0] comp1334minVal;
    wire [5:0] comp1334minI, comp1334minJ;
    Comparator comp1334(SADValues[2721*12 +: 12], 42, 33, SADValues[2784*12 +: 12], 43, 32, comp1334minVal, comp1334minI, comp1334minJ);
    wire [11:0] comp1335minVal;
    wire [5:0] comp1335minI, comp1335minJ;
    Comparator comp1335(SADValues[2847*12 +: 12], 44, 31, SADValues[2910*12 +: 12], 45, 30, comp1335minVal, comp1335minI, comp1335minJ);
    wire [11:0] comp1336minVal;
    wire [5:0] comp1336minI, comp1336minJ;
    Comparator comp1336(SADValues[2973*12 +: 12], 46, 29, SADValues[3036*12 +: 12], 47, 28, comp1336minVal, comp1336minI, comp1336minJ);
    wire [11:0] comp1337minVal;
    wire [5:0] comp1337minI, comp1337minJ;
    Comparator comp1337(SADValues[3099*12 +: 12], 48, 27, SADValues[3162*12 +: 12], 49, 26, comp1337minVal, comp1337minI, comp1337minJ);
    wire [11:0] comp1338minVal;
    wire [5:0] comp1338minI, comp1338minJ;
    Comparator comp1338(SADValues[3225*12 +: 12], 50, 25, SADValues[3288*12 +: 12], 51, 24, comp1338minVal, comp1338minI, comp1338minJ);
    wire [11:0] comp1339minVal;
    wire [5:0] comp1339minI, comp1339minJ;
    Comparator comp1339(SADValues[3351*12 +: 12], 52, 23, SADValues[3414*12 +: 12], 53, 22, comp1339minVal, comp1339minI, comp1339minJ);
    wire [11:0] comp1340minVal;
    wire [5:0] comp1340minI, comp1340minJ;
    Comparator comp1340(SADValues[3477*12 +: 12], 54, 21, SADValues[3540*12 +: 12], 55, 20, comp1340minVal, comp1340minI, comp1340minJ);
    wire [11:0] comp1341minVal;
    wire [5:0] comp1341minI, comp1341minJ;
    Comparator comp1341(SADValues[3603*12 +: 12], 56, 19, SADValues[3666*12 +: 12], 57, 18, comp1341minVal, comp1341minI, comp1341minJ);
    wire [11:0] comp1342minVal;
    wire [5:0] comp1342minI, comp1342minJ;
    Comparator comp1342(SADValues[3729*12 +: 12], 58, 17, SADValues[3792*12 +: 12], 59, 16, comp1342minVal, comp1342minI, comp1342minJ);
    wire [11:0] comp1343minVal;
    wire [5:0] comp1343minI, comp1343minJ;
    Comparator comp1343(SADValues[3855*12 +: 12], 60, 15, SADValues[3856*12 +: 12], 60, 16, comp1343minVal, comp1343minI, comp1343minJ);
    wire [11:0] comp1344minVal;
    wire [5:0] comp1344minI, comp1344minJ;
    Comparator comp1344(SADValues[3793*12 +: 12], 59, 17, SADValues[3730*12 +: 12], 58, 18, comp1344minVal, comp1344minI, comp1344minJ);
    wire [11:0] comp1345minVal;
    wire [5:0] comp1345minI, comp1345minJ;
    Comparator comp1345(SADValues[3667*12 +: 12], 57, 19, SADValues[3604*12 +: 12], 56, 20, comp1345minVal, comp1345minI, comp1345minJ);
    wire [11:0] comp1346minVal;
    wire [5:0] comp1346minI, comp1346minJ;
    Comparator comp1346(SADValues[3541*12 +: 12], 55, 21, SADValues[3478*12 +: 12], 54, 22, comp1346minVal, comp1346minI, comp1346minJ);
    wire [11:0] comp1347minVal;
    wire [5:0] comp1347minI, comp1347minJ;
    Comparator comp1347(SADValues[3415*12 +: 12], 53, 23, SADValues[3352*12 +: 12], 52, 24, comp1347minVal, comp1347minI, comp1347minJ);
    wire [11:0] comp1348minVal;
    wire [5:0] comp1348minI, comp1348minJ;
    Comparator comp1348(SADValues[3289*12 +: 12], 51, 25, SADValues[3226*12 +: 12], 50, 26, comp1348minVal, comp1348minI, comp1348minJ);
    wire [11:0] comp1349minVal;
    wire [5:0] comp1349minI, comp1349minJ;
    Comparator comp1349(SADValues[3163*12 +: 12], 49, 27, SADValues[3100*12 +: 12], 48, 28, comp1349minVal, comp1349minI, comp1349minJ);
    wire [11:0] comp1350minVal;
    wire [5:0] comp1350minI, comp1350minJ;
    Comparator comp1350(SADValues[3037*12 +: 12], 47, 29, SADValues[2974*12 +: 12], 46, 30, comp1350minVal, comp1350minI, comp1350minJ);
    wire [11:0] comp1351minVal;
    wire [5:0] comp1351minI, comp1351minJ;
    Comparator comp1351(SADValues[2911*12 +: 12], 45, 31, SADValues[2848*12 +: 12], 44, 32, comp1351minVal, comp1351minI, comp1351minJ);
    wire [11:0] comp1352minVal;
    wire [5:0] comp1352minI, comp1352minJ;
    Comparator comp1352(SADValues[2785*12 +: 12], 43, 33, SADValues[2722*12 +: 12], 42, 34, comp1352minVal, comp1352minI, comp1352minJ);
    wire [11:0] comp1353minVal;
    wire [5:0] comp1353minI, comp1353minJ;
    Comparator comp1353(SADValues[2659*12 +: 12], 41, 35, SADValues[2596*12 +: 12], 40, 36, comp1353minVal, comp1353minI, comp1353minJ);
    wire [11:0] comp1354minVal;
    wire [5:0] comp1354minI, comp1354minJ;
    Comparator comp1354(SADValues[2533*12 +: 12], 39, 37, SADValues[2470*12 +: 12], 38, 38, comp1354minVal, comp1354minI, comp1354minJ);
    wire [11:0] comp1355minVal;
    wire [5:0] comp1355minI, comp1355minJ;
    Comparator comp1355(SADValues[2407*12 +: 12], 37, 39, SADValues[2344*12 +: 12], 36, 40, comp1355minVal, comp1355minI, comp1355minJ);
    wire [11:0] comp1356minVal;
    wire [5:0] comp1356minI, comp1356minJ;
    Comparator comp1356(SADValues[2281*12 +: 12], 35, 41, SADValues[2218*12 +: 12], 34, 42, comp1356minVal, comp1356minI, comp1356minJ);
    wire [11:0] comp1357minVal;
    wire [5:0] comp1357minI, comp1357minJ;
    Comparator comp1357(SADValues[2155*12 +: 12], 33, 43, SADValues[2092*12 +: 12], 32, 44, comp1357minVal, comp1357minI, comp1357minJ);
    wire [11:0] comp1358minVal;
    wire [5:0] comp1358minI, comp1358minJ;
    Comparator comp1358(SADValues[2029*12 +: 12], 31, 45, SADValues[1966*12 +: 12], 30, 46, comp1358minVal, comp1358minI, comp1358minJ);
    wire [11:0] comp1359minVal;
    wire [5:0] comp1359minI, comp1359minJ;
    Comparator comp1359(SADValues[1903*12 +: 12], 29, 47, SADValues[1840*12 +: 12], 28, 48, comp1359minVal, comp1359minI, comp1359minJ);
    wire [11:0] comp1360minVal;
    wire [5:0] comp1360minI, comp1360minJ;
    Comparator comp1360(SADValues[1777*12 +: 12], 27, 49, SADValues[1714*12 +: 12], 26, 50, comp1360minVal, comp1360minI, comp1360minJ);
    wire [11:0] comp1361minVal;
    wire [5:0] comp1361minI, comp1361minJ;
    Comparator comp1361(SADValues[1651*12 +: 12], 25, 51, SADValues[1588*12 +: 12], 24, 52, comp1361minVal, comp1361minI, comp1361minJ);
    wire [11:0] comp1362minVal;
    wire [5:0] comp1362minI, comp1362minJ;
    Comparator comp1362(SADValues[1525*12 +: 12], 23, 53, SADValues[1462*12 +: 12], 22, 54, comp1362minVal, comp1362minI, comp1362minJ);
    wire [11:0] comp1363minVal;
    wire [5:0] comp1363minI, comp1363minJ;
    Comparator comp1363(SADValues[1399*12 +: 12], 21, 55, SADValues[1336*12 +: 12], 20, 56, comp1363minVal, comp1363minI, comp1363minJ);
    wire [11:0] comp1364minVal;
    wire [5:0] comp1364minI, comp1364minJ;
    Comparator comp1364(SADValues[1273*12 +: 12], 19, 57, SADValues[1210*12 +: 12], 18, 58, comp1364minVal, comp1364minI, comp1364minJ);
    wire [11:0] comp1365minVal;
    wire [5:0] comp1365minI, comp1365minJ;
    Comparator comp1365(SADValues[1147*12 +: 12], 17, 59, SADValues[1084*12 +: 12], 16, 60, comp1365minVal, comp1365minI, comp1365minJ);
    wire [11:0] comp1366minVal;
    wire [5:0] comp1366minI, comp1366minJ;
    Comparator comp1366(SADValues[1148*12 +: 12], 17, 60, SADValues[1211*12 +: 12], 18, 59, comp1366minVal, comp1366minI, comp1366minJ);
    wire [11:0] comp1367minVal;
    wire [5:0] comp1367minI, comp1367minJ;
    Comparator comp1367(SADValues[1274*12 +: 12], 19, 58, SADValues[1337*12 +: 12], 20, 57, comp1367minVal, comp1367minI, comp1367minJ);
    wire [11:0] comp1368minVal;
    wire [5:0] comp1368minI, comp1368minJ;
    Comparator comp1368(SADValues[1400*12 +: 12], 21, 56, SADValues[1463*12 +: 12], 22, 55, comp1368minVal, comp1368minI, comp1368minJ);
    wire [11:0] comp1369minVal;
    wire [5:0] comp1369minI, comp1369minJ;
    Comparator comp1369(SADValues[1526*12 +: 12], 23, 54, SADValues[1589*12 +: 12], 24, 53, comp1369minVal, comp1369minI, comp1369minJ);
    wire [11:0] comp1370minVal;
    wire [5:0] comp1370minI, comp1370minJ;
    Comparator comp1370(SADValues[1652*12 +: 12], 25, 52, SADValues[1715*12 +: 12], 26, 51, comp1370minVal, comp1370minI, comp1370minJ);
    wire [11:0] comp1371minVal;
    wire [5:0] comp1371minI, comp1371minJ;
    Comparator comp1371(SADValues[1778*12 +: 12], 27, 50, SADValues[1841*12 +: 12], 28, 49, comp1371minVal, comp1371minI, comp1371minJ);
    wire [11:0] comp1372minVal;
    wire [5:0] comp1372minI, comp1372minJ;
    Comparator comp1372(SADValues[1904*12 +: 12], 29, 48, SADValues[1967*12 +: 12], 30, 47, comp1372minVal, comp1372minI, comp1372minJ);
    wire [11:0] comp1373minVal;
    wire [5:0] comp1373minI, comp1373minJ;
    Comparator comp1373(SADValues[2030*12 +: 12], 31, 46, SADValues[2093*12 +: 12], 32, 45, comp1373minVal, comp1373minI, comp1373minJ);
    wire [11:0] comp1374minVal;
    wire [5:0] comp1374minI, comp1374minJ;
    Comparator comp1374(SADValues[2156*12 +: 12], 33, 44, SADValues[2219*12 +: 12], 34, 43, comp1374minVal, comp1374minI, comp1374minJ);
    wire [11:0] comp1375minVal;
    wire [5:0] comp1375minI, comp1375minJ;
    Comparator comp1375(SADValues[2282*12 +: 12], 35, 42, SADValues[2345*12 +: 12], 36, 41, comp1375minVal, comp1375minI, comp1375minJ);
    wire [11:0] comp1376minVal;
    wire [5:0] comp1376minI, comp1376minJ;
    Comparator comp1376(SADValues[2408*12 +: 12], 37, 40, SADValues[2471*12 +: 12], 38, 39, comp1376minVal, comp1376minI, comp1376minJ);
    wire [11:0] comp1377minVal;
    wire [5:0] comp1377minI, comp1377minJ;
    Comparator comp1377(SADValues[2534*12 +: 12], 39, 38, SADValues[2597*12 +: 12], 40, 37, comp1377minVal, comp1377minI, comp1377minJ);
    wire [11:0] comp1378minVal;
    wire [5:0] comp1378minI, comp1378minJ;
    Comparator comp1378(SADValues[2660*12 +: 12], 41, 36, SADValues[2723*12 +: 12], 42, 35, comp1378minVal, comp1378minI, comp1378minJ);
    wire [11:0] comp1379minVal;
    wire [5:0] comp1379minI, comp1379minJ;
    Comparator comp1379(SADValues[2786*12 +: 12], 43, 34, SADValues[2849*12 +: 12], 44, 33, comp1379minVal, comp1379minI, comp1379minJ);
    wire [11:0] comp1380minVal;
    wire [5:0] comp1380minI, comp1380minJ;
    Comparator comp1380(SADValues[2912*12 +: 12], 45, 32, SADValues[2975*12 +: 12], 46, 31, comp1380minVal, comp1380minI, comp1380minJ);
    wire [11:0] comp1381minVal;
    wire [5:0] comp1381minI, comp1381minJ;
    Comparator comp1381(SADValues[3038*12 +: 12], 47, 30, SADValues[3101*12 +: 12], 48, 29, comp1381minVal, comp1381minI, comp1381minJ);
    wire [11:0] comp1382minVal;
    wire [5:0] comp1382minI, comp1382minJ;
    Comparator comp1382(SADValues[3164*12 +: 12], 49, 28, SADValues[3227*12 +: 12], 50, 27, comp1382minVal, comp1382minI, comp1382minJ);
    wire [11:0] comp1383minVal;
    wire [5:0] comp1383minI, comp1383minJ;
    Comparator comp1383(SADValues[3290*12 +: 12], 51, 26, SADValues[3353*12 +: 12], 52, 25, comp1383minVal, comp1383minI, comp1383minJ);
    wire [11:0] comp1384minVal;
    wire [5:0] comp1384minI, comp1384minJ;
    Comparator comp1384(SADValues[3416*12 +: 12], 53, 24, SADValues[3479*12 +: 12], 54, 23, comp1384minVal, comp1384minI, comp1384minJ);
    wire [11:0] comp1385minVal;
    wire [5:0] comp1385minI, comp1385minJ;
    Comparator comp1385(SADValues[3542*12 +: 12], 55, 22, SADValues[3605*12 +: 12], 56, 21, comp1385minVal, comp1385minI, comp1385minJ);
    wire [11:0] comp1386minVal;
    wire [5:0] comp1386minI, comp1386minJ;
    Comparator comp1386(SADValues[3668*12 +: 12], 57, 20, SADValues[3731*12 +: 12], 58, 19, comp1386minVal, comp1386minI, comp1386minJ);
    wire [11:0] comp1387minVal;
    wire [5:0] comp1387minI, comp1387minJ;
    Comparator comp1387(SADValues[3794*12 +: 12], 59, 18, SADValues[3857*12 +: 12], 60, 17, comp1387minVal, comp1387minI, comp1387minJ);
    wire [11:0] comp1388minVal;
    wire [5:0] comp1388minI, comp1388minJ;
    Comparator comp1388(SADValues[3858*12 +: 12], 60, 18, SADValues[3795*12 +: 12], 59, 19, comp1388minVal, comp1388minI, comp1388minJ);
    wire [11:0] comp1389minVal;
    wire [5:0] comp1389minI, comp1389minJ;
    Comparator comp1389(SADValues[3732*12 +: 12], 58, 20, SADValues[3669*12 +: 12], 57, 21, comp1389minVal, comp1389minI, comp1389minJ);
    wire [11:0] comp1390minVal;
    wire [5:0] comp1390minI, comp1390minJ;
    Comparator comp1390(SADValues[3606*12 +: 12], 56, 22, SADValues[3543*12 +: 12], 55, 23, comp1390minVal, comp1390minI, comp1390minJ);
    wire [11:0] comp1391minVal;
    wire [5:0] comp1391minI, comp1391minJ;
    Comparator comp1391(SADValues[3480*12 +: 12], 54, 24, SADValues[3417*12 +: 12], 53, 25, comp1391minVal, comp1391minI, comp1391minJ);
    wire [11:0] comp1392minVal;
    wire [5:0] comp1392minI, comp1392minJ;
    Comparator comp1392(SADValues[3354*12 +: 12], 52, 26, SADValues[3291*12 +: 12], 51, 27, comp1392minVal, comp1392minI, comp1392minJ);
    wire [11:0] comp1393minVal;
    wire [5:0] comp1393minI, comp1393minJ;
    Comparator comp1393(SADValues[3228*12 +: 12], 50, 28, SADValues[3165*12 +: 12], 49, 29, comp1393minVal, comp1393minI, comp1393minJ);
    wire [11:0] comp1394minVal;
    wire [5:0] comp1394minI, comp1394minJ;
    Comparator comp1394(SADValues[3102*12 +: 12], 48, 30, SADValues[3039*12 +: 12], 47, 31, comp1394minVal, comp1394minI, comp1394minJ);
    wire [11:0] comp1395minVal;
    wire [5:0] comp1395minI, comp1395minJ;
    Comparator comp1395(SADValues[2976*12 +: 12], 46, 32, SADValues[2913*12 +: 12], 45, 33, comp1395minVal, comp1395minI, comp1395minJ);
    wire [11:0] comp1396minVal;
    wire [5:0] comp1396minI, comp1396minJ;
    Comparator comp1396(SADValues[2850*12 +: 12], 44, 34, SADValues[2787*12 +: 12], 43, 35, comp1396minVal, comp1396minI, comp1396minJ);
    wire [11:0] comp1397minVal;
    wire [5:0] comp1397minI, comp1397minJ;
    Comparator comp1397(SADValues[2724*12 +: 12], 42, 36, SADValues[2661*12 +: 12], 41, 37, comp1397minVal, comp1397minI, comp1397minJ);
    wire [11:0] comp1398minVal;
    wire [5:0] comp1398minI, comp1398minJ;
    Comparator comp1398(SADValues[2598*12 +: 12], 40, 38, SADValues[2535*12 +: 12], 39, 39, comp1398minVal, comp1398minI, comp1398minJ);
    wire [11:0] comp1399minVal;
    wire [5:0] comp1399minI, comp1399minJ;
    Comparator comp1399(SADValues[2472*12 +: 12], 38, 40, SADValues[2409*12 +: 12], 37, 41, comp1399minVal, comp1399minI, comp1399minJ);
    wire [11:0] comp1400minVal;
    wire [5:0] comp1400minI, comp1400minJ;
    Comparator comp1400(SADValues[2346*12 +: 12], 36, 42, SADValues[2283*12 +: 12], 35, 43, comp1400minVal, comp1400minI, comp1400minJ);
    wire [11:0] comp1401minVal;
    wire [5:0] comp1401minI, comp1401minJ;
    Comparator comp1401(SADValues[2220*12 +: 12], 34, 44, SADValues[2157*12 +: 12], 33, 45, comp1401minVal, comp1401minI, comp1401minJ);
    wire [11:0] comp1402minVal;
    wire [5:0] comp1402minI, comp1402minJ;
    Comparator comp1402(SADValues[2094*12 +: 12], 32, 46, SADValues[2031*12 +: 12], 31, 47, comp1402minVal, comp1402minI, comp1402minJ);
    wire [11:0] comp1403minVal;
    wire [5:0] comp1403minI, comp1403minJ;
    Comparator comp1403(SADValues[1968*12 +: 12], 30, 48, SADValues[1905*12 +: 12], 29, 49, comp1403minVal, comp1403minI, comp1403minJ);
    wire [11:0] comp1404minVal;
    wire [5:0] comp1404minI, comp1404minJ;
    Comparator comp1404(SADValues[1842*12 +: 12], 28, 50, SADValues[1779*12 +: 12], 27, 51, comp1404minVal, comp1404minI, comp1404minJ);
    wire [11:0] comp1405minVal;
    wire [5:0] comp1405minI, comp1405minJ;
    Comparator comp1405(SADValues[1716*12 +: 12], 26, 52, SADValues[1653*12 +: 12], 25, 53, comp1405minVal, comp1405minI, comp1405minJ);
    wire [11:0] comp1406minVal;
    wire [5:0] comp1406minI, comp1406minJ;
    Comparator comp1406(SADValues[1590*12 +: 12], 24, 54, SADValues[1527*12 +: 12], 23, 55, comp1406minVal, comp1406minI, comp1406minJ);
    wire [11:0] comp1407minVal;
    wire [5:0] comp1407minI, comp1407minJ;
    Comparator comp1407(SADValues[1464*12 +: 12], 22, 56, SADValues[1401*12 +: 12], 21, 57, comp1407minVal, comp1407minI, comp1407minJ);
    wire [11:0] comp1408minVal;
    wire [5:0] comp1408minI, comp1408minJ;
    Comparator comp1408(SADValues[1338*12 +: 12], 20, 58, SADValues[1275*12 +: 12], 19, 59, comp1408minVal, comp1408minI, comp1408minJ);
    wire [11:0] comp1409minVal;
    wire [5:0] comp1409minI, comp1409minJ;
    Comparator comp1409(SADValues[1212*12 +: 12], 18, 60, SADValues[1276*12 +: 12], 19, 60, comp1409minVal, comp1409minI, comp1409minJ);
    wire [11:0] comp1410minVal;
    wire [5:0] comp1410minI, comp1410minJ;
    Comparator comp1410(SADValues[1339*12 +: 12], 20, 59, SADValues[1402*12 +: 12], 21, 58, comp1410minVal, comp1410minI, comp1410minJ);
    wire [11:0] comp1411minVal;
    wire [5:0] comp1411minI, comp1411minJ;
    Comparator comp1411(SADValues[1465*12 +: 12], 22, 57, SADValues[1528*12 +: 12], 23, 56, comp1411minVal, comp1411minI, comp1411minJ);
    wire [11:0] comp1412minVal;
    wire [5:0] comp1412minI, comp1412minJ;
    Comparator comp1412(SADValues[1591*12 +: 12], 24, 55, SADValues[1654*12 +: 12], 25, 54, comp1412minVal, comp1412minI, comp1412minJ);
    wire [11:0] comp1413minVal;
    wire [5:0] comp1413minI, comp1413minJ;
    Comparator comp1413(SADValues[1717*12 +: 12], 26, 53, SADValues[1780*12 +: 12], 27, 52, comp1413minVal, comp1413minI, comp1413minJ);
    wire [11:0] comp1414minVal;
    wire [5:0] comp1414minI, comp1414minJ;
    Comparator comp1414(SADValues[1843*12 +: 12], 28, 51, SADValues[1906*12 +: 12], 29, 50, comp1414minVal, comp1414minI, comp1414minJ);
    wire [11:0] comp1415minVal;
    wire [5:0] comp1415minI, comp1415minJ;
    Comparator comp1415(SADValues[1969*12 +: 12], 30, 49, SADValues[2032*12 +: 12], 31, 48, comp1415minVal, comp1415minI, comp1415minJ);
    wire [11:0] comp1416minVal;
    wire [5:0] comp1416minI, comp1416minJ;
    Comparator comp1416(SADValues[2095*12 +: 12], 32, 47, SADValues[2158*12 +: 12], 33, 46, comp1416minVal, comp1416minI, comp1416minJ);
    wire [11:0] comp1417minVal;
    wire [5:0] comp1417minI, comp1417minJ;
    Comparator comp1417(SADValues[2221*12 +: 12], 34, 45, SADValues[2284*12 +: 12], 35, 44, comp1417minVal, comp1417minI, comp1417minJ);
    wire [11:0] comp1418minVal;
    wire [5:0] comp1418minI, comp1418minJ;
    Comparator comp1418(SADValues[2347*12 +: 12], 36, 43, SADValues[2410*12 +: 12], 37, 42, comp1418minVal, comp1418minI, comp1418minJ);
    wire [11:0] comp1419minVal;
    wire [5:0] comp1419minI, comp1419minJ;
    Comparator comp1419(SADValues[2473*12 +: 12], 38, 41, SADValues[2536*12 +: 12], 39, 40, comp1419minVal, comp1419minI, comp1419minJ);
    wire [11:0] comp1420minVal;
    wire [5:0] comp1420minI, comp1420minJ;
    Comparator comp1420(SADValues[2599*12 +: 12], 40, 39, SADValues[2662*12 +: 12], 41, 38, comp1420minVal, comp1420minI, comp1420minJ);
    wire [11:0] comp1421minVal;
    wire [5:0] comp1421minI, comp1421minJ;
    Comparator comp1421(SADValues[2725*12 +: 12], 42, 37, SADValues[2788*12 +: 12], 43, 36, comp1421minVal, comp1421minI, comp1421minJ);
    wire [11:0] comp1422minVal;
    wire [5:0] comp1422minI, comp1422minJ;
    Comparator comp1422(SADValues[2851*12 +: 12], 44, 35, SADValues[2914*12 +: 12], 45, 34, comp1422minVal, comp1422minI, comp1422minJ);
    wire [11:0] comp1423minVal;
    wire [5:0] comp1423minI, comp1423minJ;
    Comparator comp1423(SADValues[2977*12 +: 12], 46, 33, SADValues[3040*12 +: 12], 47, 32, comp1423minVal, comp1423minI, comp1423minJ);
    wire [11:0] comp1424minVal;
    wire [5:0] comp1424minI, comp1424minJ;
    Comparator comp1424(SADValues[3103*12 +: 12], 48, 31, SADValues[3166*12 +: 12], 49, 30, comp1424minVal, comp1424minI, comp1424minJ);
    wire [11:0] comp1425minVal;
    wire [5:0] comp1425minI, comp1425minJ;
    Comparator comp1425(SADValues[3229*12 +: 12], 50, 29, SADValues[3292*12 +: 12], 51, 28, comp1425minVal, comp1425minI, comp1425minJ);
    wire [11:0] comp1426minVal;
    wire [5:0] comp1426minI, comp1426minJ;
    Comparator comp1426(SADValues[3355*12 +: 12], 52, 27, SADValues[3418*12 +: 12], 53, 26, comp1426minVal, comp1426minI, comp1426minJ);
    wire [11:0] comp1427minVal;
    wire [5:0] comp1427minI, comp1427minJ;
    Comparator comp1427(SADValues[3481*12 +: 12], 54, 25, SADValues[3544*12 +: 12], 55, 24, comp1427minVal, comp1427minI, comp1427minJ);
    wire [11:0] comp1428minVal;
    wire [5:0] comp1428minI, comp1428minJ;
    Comparator comp1428(SADValues[3607*12 +: 12], 56, 23, SADValues[3670*12 +: 12], 57, 22, comp1428minVal, comp1428minI, comp1428minJ);
    wire [11:0] comp1429minVal;
    wire [5:0] comp1429minI, comp1429minJ;
    Comparator comp1429(SADValues[3733*12 +: 12], 58, 21, SADValues[3796*12 +: 12], 59, 20, comp1429minVal, comp1429minI, comp1429minJ);
    wire [11:0] comp1430minVal;
    wire [5:0] comp1430minI, comp1430minJ;
    Comparator comp1430(SADValues[3859*12 +: 12], 60, 19, SADValues[3860*12 +: 12], 60, 20, comp1430minVal, comp1430minI, comp1430minJ);
    wire [11:0] comp1431minVal;
    wire [5:0] comp1431minI, comp1431minJ;
    Comparator comp1431(SADValues[3797*12 +: 12], 59, 21, SADValues[3734*12 +: 12], 58, 22, comp1431minVal, comp1431minI, comp1431minJ);
    wire [11:0] comp1432minVal;
    wire [5:0] comp1432minI, comp1432minJ;
    Comparator comp1432(SADValues[3671*12 +: 12], 57, 23, SADValues[3608*12 +: 12], 56, 24, comp1432minVal, comp1432minI, comp1432minJ);
    wire [11:0] comp1433minVal;
    wire [5:0] comp1433minI, comp1433minJ;
    Comparator comp1433(SADValues[3545*12 +: 12], 55, 25, SADValues[3482*12 +: 12], 54, 26, comp1433minVal, comp1433minI, comp1433minJ);
    wire [11:0] comp1434minVal;
    wire [5:0] comp1434minI, comp1434minJ;
    Comparator comp1434(SADValues[3419*12 +: 12], 53, 27, SADValues[3356*12 +: 12], 52, 28, comp1434minVal, comp1434minI, comp1434minJ);
    wire [11:0] comp1435minVal;
    wire [5:0] comp1435minI, comp1435minJ;
    Comparator comp1435(SADValues[3293*12 +: 12], 51, 29, SADValues[3230*12 +: 12], 50, 30, comp1435minVal, comp1435minI, comp1435minJ);
    wire [11:0] comp1436minVal;
    wire [5:0] comp1436minI, comp1436minJ;
    Comparator comp1436(SADValues[3167*12 +: 12], 49, 31, SADValues[3104*12 +: 12], 48, 32, comp1436minVal, comp1436minI, comp1436minJ);
    wire [11:0] comp1437minVal;
    wire [5:0] comp1437minI, comp1437minJ;
    Comparator comp1437(SADValues[3041*12 +: 12], 47, 33, SADValues[2978*12 +: 12], 46, 34, comp1437minVal, comp1437minI, comp1437minJ);
    wire [11:0] comp1438minVal;
    wire [5:0] comp1438minI, comp1438minJ;
    Comparator comp1438(SADValues[2915*12 +: 12], 45, 35, SADValues[2852*12 +: 12], 44, 36, comp1438minVal, comp1438minI, comp1438minJ);
    wire [11:0] comp1439minVal;
    wire [5:0] comp1439minI, comp1439minJ;
    Comparator comp1439(SADValues[2789*12 +: 12], 43, 37, SADValues[2726*12 +: 12], 42, 38, comp1439minVal, comp1439minI, comp1439minJ);
    wire [11:0] comp1440minVal;
    wire [5:0] comp1440minI, comp1440minJ;
    Comparator comp1440(SADValues[2663*12 +: 12], 41, 39, SADValues[2600*12 +: 12], 40, 40, comp1440minVal, comp1440minI, comp1440minJ);
    wire [11:0] comp1441minVal;
    wire [5:0] comp1441minI, comp1441minJ;
    Comparator comp1441(SADValues[2537*12 +: 12], 39, 41, SADValues[2474*12 +: 12], 38, 42, comp1441minVal, comp1441minI, comp1441minJ);
    wire [11:0] comp1442minVal;
    wire [5:0] comp1442minI, comp1442minJ;
    Comparator comp1442(SADValues[2411*12 +: 12], 37, 43, SADValues[2348*12 +: 12], 36, 44, comp1442minVal, comp1442minI, comp1442minJ);
    wire [11:0] comp1443minVal;
    wire [5:0] comp1443minI, comp1443minJ;
    Comparator comp1443(SADValues[2285*12 +: 12], 35, 45, SADValues[2222*12 +: 12], 34, 46, comp1443minVal, comp1443minI, comp1443minJ);
    wire [11:0] comp1444minVal;
    wire [5:0] comp1444minI, comp1444minJ;
    Comparator comp1444(SADValues[2159*12 +: 12], 33, 47, SADValues[2096*12 +: 12], 32, 48, comp1444minVal, comp1444minI, comp1444minJ);
    wire [11:0] comp1445minVal;
    wire [5:0] comp1445minI, comp1445minJ;
    Comparator comp1445(SADValues[2033*12 +: 12], 31, 49, SADValues[1970*12 +: 12], 30, 50, comp1445minVal, comp1445minI, comp1445minJ);
    wire [11:0] comp1446minVal;
    wire [5:0] comp1446minI, comp1446minJ;
    Comparator comp1446(SADValues[1907*12 +: 12], 29, 51, SADValues[1844*12 +: 12], 28, 52, comp1446minVal, comp1446minI, comp1446minJ);
    wire [11:0] comp1447minVal;
    wire [5:0] comp1447minI, comp1447minJ;
    Comparator comp1447(SADValues[1781*12 +: 12], 27, 53, SADValues[1718*12 +: 12], 26, 54, comp1447minVal, comp1447minI, comp1447minJ);
    wire [11:0] comp1448minVal;
    wire [5:0] comp1448minI, comp1448minJ;
    Comparator comp1448(SADValues[1655*12 +: 12], 25, 55, SADValues[1592*12 +: 12], 24, 56, comp1448minVal, comp1448minI, comp1448minJ);
    wire [11:0] comp1449minVal;
    wire [5:0] comp1449minI, comp1449minJ;
    Comparator comp1449(SADValues[1529*12 +: 12], 23, 57, SADValues[1466*12 +: 12], 22, 58, comp1449minVal, comp1449minI, comp1449minJ);
    wire [11:0] comp1450minVal;
    wire [5:0] comp1450minI, comp1450minJ;
    Comparator comp1450(SADValues[1403*12 +: 12], 21, 59, SADValues[1340*12 +: 12], 20, 60, comp1450minVal, comp1450minI, comp1450minJ);
    wire [11:0] comp1451minVal;
    wire [5:0] comp1451minI, comp1451minJ;
    Comparator comp1451(SADValues[1404*12 +: 12], 21, 60, SADValues[1467*12 +: 12], 22, 59, comp1451minVal, comp1451minI, comp1451minJ);
    wire [11:0] comp1452minVal;
    wire [5:0] comp1452minI, comp1452minJ;
    Comparator comp1452(SADValues[1530*12 +: 12], 23, 58, SADValues[1593*12 +: 12], 24, 57, comp1452minVal, comp1452minI, comp1452minJ);
    wire [11:0] comp1453minVal;
    wire [5:0] comp1453minI, comp1453minJ;
    Comparator comp1453(SADValues[1656*12 +: 12], 25, 56, SADValues[1719*12 +: 12], 26, 55, comp1453minVal, comp1453minI, comp1453minJ);
    wire [11:0] comp1454minVal;
    wire [5:0] comp1454minI, comp1454minJ;
    Comparator comp1454(SADValues[1782*12 +: 12], 27, 54, SADValues[1845*12 +: 12], 28, 53, comp1454minVal, comp1454minI, comp1454minJ);
    wire [11:0] comp1455minVal;
    wire [5:0] comp1455minI, comp1455minJ;
    Comparator comp1455(SADValues[1908*12 +: 12], 29, 52, SADValues[1971*12 +: 12], 30, 51, comp1455minVal, comp1455minI, comp1455minJ);
    wire [11:0] comp1456minVal;
    wire [5:0] comp1456minI, comp1456minJ;
    Comparator comp1456(SADValues[2034*12 +: 12], 31, 50, SADValues[2097*12 +: 12], 32, 49, comp1456minVal, comp1456minI, comp1456minJ);
    wire [11:0] comp1457minVal;
    wire [5:0] comp1457minI, comp1457minJ;
    Comparator comp1457(SADValues[2160*12 +: 12], 33, 48, SADValues[2223*12 +: 12], 34, 47, comp1457minVal, comp1457minI, comp1457minJ);
    wire [11:0] comp1458minVal;
    wire [5:0] comp1458minI, comp1458minJ;
    Comparator comp1458(SADValues[2286*12 +: 12], 35, 46, SADValues[2349*12 +: 12], 36, 45, comp1458minVal, comp1458minI, comp1458minJ);
    wire [11:0] comp1459minVal;
    wire [5:0] comp1459minI, comp1459minJ;
    Comparator comp1459(SADValues[2412*12 +: 12], 37, 44, SADValues[2475*12 +: 12], 38, 43, comp1459minVal, comp1459minI, comp1459minJ);
    wire [11:0] comp1460minVal;
    wire [5:0] comp1460minI, comp1460minJ;
    Comparator comp1460(SADValues[2538*12 +: 12], 39, 42, SADValues[2601*12 +: 12], 40, 41, comp1460minVal, comp1460minI, comp1460minJ);
    wire [11:0] comp1461minVal;
    wire [5:0] comp1461minI, comp1461minJ;
    Comparator comp1461(SADValues[2664*12 +: 12], 41, 40, SADValues[2727*12 +: 12], 42, 39, comp1461minVal, comp1461minI, comp1461minJ);
    wire [11:0] comp1462minVal;
    wire [5:0] comp1462minI, comp1462minJ;
    Comparator comp1462(SADValues[2790*12 +: 12], 43, 38, SADValues[2853*12 +: 12], 44, 37, comp1462minVal, comp1462minI, comp1462minJ);
    wire [11:0] comp1463minVal;
    wire [5:0] comp1463minI, comp1463minJ;
    Comparator comp1463(SADValues[2916*12 +: 12], 45, 36, SADValues[2979*12 +: 12], 46, 35, comp1463minVal, comp1463minI, comp1463minJ);
    wire [11:0] comp1464minVal;
    wire [5:0] comp1464minI, comp1464minJ;
    Comparator comp1464(SADValues[3042*12 +: 12], 47, 34, SADValues[3105*12 +: 12], 48, 33, comp1464minVal, comp1464minI, comp1464minJ);
    wire [11:0] comp1465minVal;
    wire [5:0] comp1465minI, comp1465minJ;
    Comparator comp1465(SADValues[3168*12 +: 12], 49, 32, SADValues[3231*12 +: 12], 50, 31, comp1465minVal, comp1465minI, comp1465minJ);
    wire [11:0] comp1466minVal;
    wire [5:0] comp1466minI, comp1466minJ;
    Comparator comp1466(SADValues[3294*12 +: 12], 51, 30, SADValues[3357*12 +: 12], 52, 29, comp1466minVal, comp1466minI, comp1466minJ);
    wire [11:0] comp1467minVal;
    wire [5:0] comp1467minI, comp1467minJ;
    Comparator comp1467(SADValues[3420*12 +: 12], 53, 28, SADValues[3483*12 +: 12], 54, 27, comp1467minVal, comp1467minI, comp1467minJ);
    wire [11:0] comp1468minVal;
    wire [5:0] comp1468minI, comp1468minJ;
    Comparator comp1468(SADValues[3546*12 +: 12], 55, 26, SADValues[3609*12 +: 12], 56, 25, comp1468minVal, comp1468minI, comp1468minJ);
    wire [11:0] comp1469minVal;
    wire [5:0] comp1469minI, comp1469minJ;
    Comparator comp1469(SADValues[3672*12 +: 12], 57, 24, SADValues[3735*12 +: 12], 58, 23, comp1469minVal, comp1469minI, comp1469minJ);
    wire [11:0] comp1470minVal;
    wire [5:0] comp1470minI, comp1470minJ;
    Comparator comp1470(SADValues[3798*12 +: 12], 59, 22, SADValues[3861*12 +: 12], 60, 21, comp1470minVal, comp1470minI, comp1470minJ);
    wire [11:0] comp1471minVal;
    wire [5:0] comp1471minI, comp1471minJ;
    Comparator comp1471(SADValues[3862*12 +: 12], 60, 22, SADValues[3799*12 +: 12], 59, 23, comp1471minVal, comp1471minI, comp1471minJ);
    wire [11:0] comp1472minVal;
    wire [5:0] comp1472minI, comp1472minJ;
    Comparator comp1472(SADValues[3736*12 +: 12], 58, 24, SADValues[3673*12 +: 12], 57, 25, comp1472minVal, comp1472minI, comp1472minJ);
    wire [11:0] comp1473minVal;
    wire [5:0] comp1473minI, comp1473minJ;
    Comparator comp1473(SADValues[3610*12 +: 12], 56, 26, SADValues[3547*12 +: 12], 55, 27, comp1473minVal, comp1473minI, comp1473minJ);
    wire [11:0] comp1474minVal;
    wire [5:0] comp1474minI, comp1474minJ;
    Comparator comp1474(SADValues[3484*12 +: 12], 54, 28, SADValues[3421*12 +: 12], 53, 29, comp1474minVal, comp1474minI, comp1474minJ);
    wire [11:0] comp1475minVal;
    wire [5:0] comp1475minI, comp1475minJ;
    Comparator comp1475(SADValues[3358*12 +: 12], 52, 30, SADValues[3295*12 +: 12], 51, 31, comp1475minVal, comp1475minI, comp1475minJ);
    wire [11:0] comp1476minVal;
    wire [5:0] comp1476minI, comp1476minJ;
    Comparator comp1476(SADValues[3232*12 +: 12], 50, 32, SADValues[3169*12 +: 12], 49, 33, comp1476minVal, comp1476minI, comp1476minJ);
    wire [11:0] comp1477minVal;
    wire [5:0] comp1477minI, comp1477minJ;
    Comparator comp1477(SADValues[3106*12 +: 12], 48, 34, SADValues[3043*12 +: 12], 47, 35, comp1477minVal, comp1477minI, comp1477minJ);
    wire [11:0] comp1478minVal;
    wire [5:0] comp1478minI, comp1478minJ;
    Comparator comp1478(SADValues[2980*12 +: 12], 46, 36, SADValues[2917*12 +: 12], 45, 37, comp1478minVal, comp1478minI, comp1478minJ);
    wire [11:0] comp1479minVal;
    wire [5:0] comp1479minI, comp1479minJ;
    Comparator comp1479(SADValues[2854*12 +: 12], 44, 38, SADValues[2791*12 +: 12], 43, 39, comp1479minVal, comp1479minI, comp1479minJ);
    wire [11:0] comp1480minVal;
    wire [5:0] comp1480minI, comp1480minJ;
    Comparator comp1480(SADValues[2728*12 +: 12], 42, 40, SADValues[2665*12 +: 12], 41, 41, comp1480minVal, comp1480minI, comp1480minJ);
    wire [11:0] comp1481minVal;
    wire [5:0] comp1481minI, comp1481minJ;
    Comparator comp1481(SADValues[2602*12 +: 12], 40, 42, SADValues[2539*12 +: 12], 39, 43, comp1481minVal, comp1481minI, comp1481minJ);
    wire [11:0] comp1482minVal;
    wire [5:0] comp1482minI, comp1482minJ;
    Comparator comp1482(SADValues[2476*12 +: 12], 38, 44, SADValues[2413*12 +: 12], 37, 45, comp1482minVal, comp1482minI, comp1482minJ);
    wire [11:0] comp1483minVal;
    wire [5:0] comp1483minI, comp1483minJ;
    Comparator comp1483(SADValues[2350*12 +: 12], 36, 46, SADValues[2287*12 +: 12], 35, 47, comp1483minVal, comp1483minI, comp1483minJ);
    wire [11:0] comp1484minVal;
    wire [5:0] comp1484minI, comp1484minJ;
    Comparator comp1484(SADValues[2224*12 +: 12], 34, 48, SADValues[2161*12 +: 12], 33, 49, comp1484minVal, comp1484minI, comp1484minJ);
    wire [11:0] comp1485minVal;
    wire [5:0] comp1485minI, comp1485minJ;
    Comparator comp1485(SADValues[2098*12 +: 12], 32, 50, SADValues[2035*12 +: 12], 31, 51, comp1485minVal, comp1485minI, comp1485minJ);
    wire [11:0] comp1486minVal;
    wire [5:0] comp1486minI, comp1486minJ;
    Comparator comp1486(SADValues[1972*12 +: 12], 30, 52, SADValues[1909*12 +: 12], 29, 53, comp1486minVal, comp1486minI, comp1486minJ);
    wire [11:0] comp1487minVal;
    wire [5:0] comp1487minI, comp1487minJ;
    Comparator comp1487(SADValues[1846*12 +: 12], 28, 54, SADValues[1783*12 +: 12], 27, 55, comp1487minVal, comp1487minI, comp1487minJ);
    wire [11:0] comp1488minVal;
    wire [5:0] comp1488minI, comp1488minJ;
    Comparator comp1488(SADValues[1720*12 +: 12], 26, 56, SADValues[1657*12 +: 12], 25, 57, comp1488minVal, comp1488minI, comp1488minJ);
    wire [11:0] comp1489minVal;
    wire [5:0] comp1489minI, comp1489minJ;
    Comparator comp1489(SADValues[1594*12 +: 12], 24, 58, SADValues[1531*12 +: 12], 23, 59, comp1489minVal, comp1489minI, comp1489minJ);
    wire [11:0] comp1490minVal;
    wire [5:0] comp1490minI, comp1490minJ;
    Comparator comp1490(SADValues[1468*12 +: 12], 22, 60, SADValues[1532*12 +: 12], 23, 60, comp1490minVal, comp1490minI, comp1490minJ);
    wire [11:0] comp1491minVal;
    wire [5:0] comp1491minI, comp1491minJ;
    Comparator comp1491(SADValues[1595*12 +: 12], 24, 59, SADValues[1658*12 +: 12], 25, 58, comp1491minVal, comp1491minI, comp1491minJ);
    wire [11:0] comp1492minVal;
    wire [5:0] comp1492minI, comp1492minJ;
    Comparator comp1492(SADValues[1721*12 +: 12], 26, 57, SADValues[1784*12 +: 12], 27, 56, comp1492minVal, comp1492minI, comp1492minJ);
    wire [11:0] comp1493minVal;
    wire [5:0] comp1493minI, comp1493minJ;
    Comparator comp1493(SADValues[1847*12 +: 12], 28, 55, SADValues[1910*12 +: 12], 29, 54, comp1493minVal, comp1493minI, comp1493minJ);
    wire [11:0] comp1494minVal;
    wire [5:0] comp1494minI, comp1494minJ;
    Comparator comp1494(SADValues[1973*12 +: 12], 30, 53, SADValues[2036*12 +: 12], 31, 52, comp1494minVal, comp1494minI, comp1494minJ);
    wire [11:0] comp1495minVal;
    wire [5:0] comp1495minI, comp1495minJ;
    Comparator comp1495(SADValues[2099*12 +: 12], 32, 51, SADValues[2162*12 +: 12], 33, 50, comp1495minVal, comp1495minI, comp1495minJ);
    wire [11:0] comp1496minVal;
    wire [5:0] comp1496minI, comp1496minJ;
    Comparator comp1496(SADValues[2225*12 +: 12], 34, 49, SADValues[2288*12 +: 12], 35, 48, comp1496minVal, comp1496minI, comp1496minJ);
    wire [11:0] comp1497minVal;
    wire [5:0] comp1497minI, comp1497minJ;
    Comparator comp1497(SADValues[2351*12 +: 12], 36, 47, SADValues[2414*12 +: 12], 37, 46, comp1497minVal, comp1497minI, comp1497minJ);
    wire [11:0] comp1498minVal;
    wire [5:0] comp1498minI, comp1498minJ;
    Comparator comp1498(SADValues[2477*12 +: 12], 38, 45, SADValues[2540*12 +: 12], 39, 44, comp1498minVal, comp1498minI, comp1498minJ);
    wire [11:0] comp1499minVal;
    wire [5:0] comp1499minI, comp1499minJ;
    Comparator comp1499(SADValues[2603*12 +: 12], 40, 43, SADValues[2666*12 +: 12], 41, 42, comp1499minVal, comp1499minI, comp1499minJ);
    wire [11:0] comp1500minVal;
    wire [5:0] comp1500minI, comp1500minJ;
    Comparator comp1500(SADValues[2729*12 +: 12], 42, 41, SADValues[2792*12 +: 12], 43, 40, comp1500minVal, comp1500minI, comp1500minJ);
    wire [11:0] comp1501minVal;
    wire [5:0] comp1501minI, comp1501minJ;
    Comparator comp1501(SADValues[2855*12 +: 12], 44, 39, SADValues[2918*12 +: 12], 45, 38, comp1501minVal, comp1501minI, comp1501minJ);
    wire [11:0] comp1502minVal;
    wire [5:0] comp1502minI, comp1502minJ;
    Comparator comp1502(SADValues[2981*12 +: 12], 46, 37, SADValues[3044*12 +: 12], 47, 36, comp1502minVal, comp1502minI, comp1502minJ);
    wire [11:0] comp1503minVal;
    wire [5:0] comp1503minI, comp1503minJ;
    Comparator comp1503(SADValues[3107*12 +: 12], 48, 35, SADValues[3170*12 +: 12], 49, 34, comp1503minVal, comp1503minI, comp1503minJ);
    wire [11:0] comp1504minVal;
    wire [5:0] comp1504minI, comp1504minJ;
    Comparator comp1504(SADValues[3233*12 +: 12], 50, 33, SADValues[3296*12 +: 12], 51, 32, comp1504minVal, comp1504minI, comp1504minJ);
    wire [11:0] comp1505minVal;
    wire [5:0] comp1505minI, comp1505minJ;
    Comparator comp1505(SADValues[3359*12 +: 12], 52, 31, SADValues[3422*12 +: 12], 53, 30, comp1505minVal, comp1505minI, comp1505minJ);
    wire [11:0] comp1506minVal;
    wire [5:0] comp1506minI, comp1506minJ;
    Comparator comp1506(SADValues[3485*12 +: 12], 54, 29, SADValues[3548*12 +: 12], 55, 28, comp1506minVal, comp1506minI, comp1506minJ);
    wire [11:0] comp1507minVal;
    wire [5:0] comp1507minI, comp1507minJ;
    Comparator comp1507(SADValues[3611*12 +: 12], 56, 27, SADValues[3674*12 +: 12], 57, 26, comp1507minVal, comp1507minI, comp1507minJ);
    wire [11:0] comp1508minVal;
    wire [5:0] comp1508minI, comp1508minJ;
    Comparator comp1508(SADValues[3737*12 +: 12], 58, 25, SADValues[3800*12 +: 12], 59, 24, comp1508minVal, comp1508minI, comp1508minJ);
    wire [11:0] comp1509minVal;
    wire [5:0] comp1509minI, comp1509minJ;
    Comparator comp1509(SADValues[3863*12 +: 12], 60, 23, SADValues[3864*12 +: 12], 60, 24, comp1509minVal, comp1509minI, comp1509minJ);
    wire [11:0] comp1510minVal;
    wire [5:0] comp1510minI, comp1510minJ;
    Comparator comp1510(SADValues[3801*12 +: 12], 59, 25, SADValues[3738*12 +: 12], 58, 26, comp1510minVal, comp1510minI, comp1510minJ);
    wire [11:0] comp1511minVal;
    wire [5:0] comp1511minI, comp1511minJ;
    Comparator comp1511(SADValues[3675*12 +: 12], 57, 27, SADValues[3612*12 +: 12], 56, 28, comp1511minVal, comp1511minI, comp1511minJ);
    wire [11:0] comp1512minVal;
    wire [5:0] comp1512minI, comp1512minJ;
    Comparator comp1512(SADValues[3549*12 +: 12], 55, 29, SADValues[3486*12 +: 12], 54, 30, comp1512minVal, comp1512minI, comp1512minJ);
    wire [11:0] comp1513minVal;
    wire [5:0] comp1513minI, comp1513minJ;
    Comparator comp1513(SADValues[3423*12 +: 12], 53, 31, SADValues[3360*12 +: 12], 52, 32, comp1513minVal, comp1513minI, comp1513minJ);
    wire [11:0] comp1514minVal;
    wire [5:0] comp1514minI, comp1514minJ;
    Comparator comp1514(SADValues[3297*12 +: 12], 51, 33, SADValues[3234*12 +: 12], 50, 34, comp1514minVal, comp1514minI, comp1514minJ);
    wire [11:0] comp1515minVal;
    wire [5:0] comp1515minI, comp1515minJ;
    Comparator comp1515(SADValues[3171*12 +: 12], 49, 35, SADValues[3108*12 +: 12], 48, 36, comp1515minVal, comp1515minI, comp1515minJ);
    wire [11:0] comp1516minVal;
    wire [5:0] comp1516minI, comp1516minJ;
    Comparator comp1516(SADValues[3045*12 +: 12], 47, 37, SADValues[2982*12 +: 12], 46, 38, comp1516minVal, comp1516minI, comp1516minJ);
    wire [11:0] comp1517minVal;
    wire [5:0] comp1517minI, comp1517minJ;
    Comparator comp1517(SADValues[2919*12 +: 12], 45, 39, SADValues[2856*12 +: 12], 44, 40, comp1517minVal, comp1517minI, comp1517minJ);
    wire [11:0] comp1518minVal;
    wire [5:0] comp1518minI, comp1518minJ;
    Comparator comp1518(SADValues[2793*12 +: 12], 43, 41, SADValues[2730*12 +: 12], 42, 42, comp1518minVal, comp1518minI, comp1518minJ);
    wire [11:0] comp1519minVal;
    wire [5:0] comp1519minI, comp1519minJ;
    Comparator comp1519(SADValues[2667*12 +: 12], 41, 43, SADValues[2604*12 +: 12], 40, 44, comp1519minVal, comp1519minI, comp1519minJ);
    wire [11:0] comp1520minVal;
    wire [5:0] comp1520minI, comp1520minJ;
    Comparator comp1520(SADValues[2541*12 +: 12], 39, 45, SADValues[2478*12 +: 12], 38, 46, comp1520minVal, comp1520minI, comp1520minJ);
    wire [11:0] comp1521minVal;
    wire [5:0] comp1521minI, comp1521minJ;
    Comparator comp1521(SADValues[2415*12 +: 12], 37, 47, SADValues[2352*12 +: 12], 36, 48, comp1521minVal, comp1521minI, comp1521minJ);
    wire [11:0] comp1522minVal;
    wire [5:0] comp1522minI, comp1522minJ;
    Comparator comp1522(SADValues[2289*12 +: 12], 35, 49, SADValues[2226*12 +: 12], 34, 50, comp1522minVal, comp1522minI, comp1522minJ);
    wire [11:0] comp1523minVal;
    wire [5:0] comp1523minI, comp1523minJ;
    Comparator comp1523(SADValues[2163*12 +: 12], 33, 51, SADValues[2100*12 +: 12], 32, 52, comp1523minVal, comp1523minI, comp1523minJ);
    wire [11:0] comp1524minVal;
    wire [5:0] comp1524minI, comp1524minJ;
    Comparator comp1524(SADValues[2037*12 +: 12], 31, 53, SADValues[1974*12 +: 12], 30, 54, comp1524minVal, comp1524minI, comp1524minJ);
    wire [11:0] comp1525minVal;
    wire [5:0] comp1525minI, comp1525minJ;
    Comparator comp1525(SADValues[1911*12 +: 12], 29, 55, SADValues[1848*12 +: 12], 28, 56, comp1525minVal, comp1525minI, comp1525minJ);
    wire [11:0] comp1526minVal;
    wire [5:0] comp1526minI, comp1526minJ;
    Comparator comp1526(SADValues[1785*12 +: 12], 27, 57, SADValues[1722*12 +: 12], 26, 58, comp1526minVal, comp1526minI, comp1526minJ);
    wire [11:0] comp1527minVal;
    wire [5:0] comp1527minI, comp1527minJ;
    Comparator comp1527(SADValues[1659*12 +: 12], 25, 59, SADValues[1596*12 +: 12], 24, 60, comp1527minVal, comp1527minI, comp1527minJ);
    wire [11:0] comp1528minVal;
    wire [5:0] comp1528minI, comp1528minJ;
    Comparator comp1528(SADValues[1660*12 +: 12], 25, 60, SADValues[1723*12 +: 12], 26, 59, comp1528minVal, comp1528minI, comp1528minJ);
    wire [11:0] comp1529minVal;
    wire [5:0] comp1529minI, comp1529minJ;
    Comparator comp1529(SADValues[1786*12 +: 12], 27, 58, SADValues[1849*12 +: 12], 28, 57, comp1529minVal, comp1529minI, comp1529minJ);
    wire [11:0] comp1530minVal;
    wire [5:0] comp1530minI, comp1530minJ;
    Comparator comp1530(SADValues[1912*12 +: 12], 29, 56, SADValues[1975*12 +: 12], 30, 55, comp1530minVal, comp1530minI, comp1530minJ);
    wire [11:0] comp1531minVal;
    wire [5:0] comp1531minI, comp1531minJ;
    Comparator comp1531(SADValues[2038*12 +: 12], 31, 54, SADValues[2101*12 +: 12], 32, 53, comp1531minVal, comp1531minI, comp1531minJ);
    wire [11:0] comp1532minVal;
    wire [5:0] comp1532minI, comp1532minJ;
    Comparator comp1532(SADValues[2164*12 +: 12], 33, 52, SADValues[2227*12 +: 12], 34, 51, comp1532minVal, comp1532minI, comp1532minJ);
    wire [11:0] comp1533minVal;
    wire [5:0] comp1533minI, comp1533minJ;
    Comparator comp1533(SADValues[2290*12 +: 12], 35, 50, SADValues[2353*12 +: 12], 36, 49, comp1533minVal, comp1533minI, comp1533minJ);
    wire [11:0] comp1534minVal;
    wire [5:0] comp1534minI, comp1534minJ;
    Comparator comp1534(SADValues[2416*12 +: 12], 37, 48, SADValues[2479*12 +: 12], 38, 47, comp1534minVal, comp1534minI, comp1534minJ);
    wire [11:0] comp1535minVal;
    wire [5:0] comp1535minI, comp1535minJ;
    Comparator comp1535(SADValues[2542*12 +: 12], 39, 46, SADValues[2605*12 +: 12], 40, 45, comp1535minVal, comp1535minI, comp1535minJ);
    wire [11:0] comp1536minVal;
    wire [5:0] comp1536minI, comp1536minJ;
    Comparator comp1536(SADValues[2668*12 +: 12], 41, 44, SADValues[2731*12 +: 12], 42, 43, comp1536minVal, comp1536minI, comp1536minJ);
    wire [11:0] comp1537minVal;
    wire [5:0] comp1537minI, comp1537minJ;
    Comparator comp1537(SADValues[2794*12 +: 12], 43, 42, SADValues[2857*12 +: 12], 44, 41, comp1537minVal, comp1537minI, comp1537minJ);
    wire [11:0] comp1538minVal;
    wire [5:0] comp1538minI, comp1538minJ;
    Comparator comp1538(SADValues[2920*12 +: 12], 45, 40, SADValues[2983*12 +: 12], 46, 39, comp1538minVal, comp1538minI, comp1538minJ);
    wire [11:0] comp1539minVal;
    wire [5:0] comp1539minI, comp1539minJ;
    Comparator comp1539(SADValues[3046*12 +: 12], 47, 38, SADValues[3109*12 +: 12], 48, 37, comp1539minVal, comp1539minI, comp1539minJ);
    wire [11:0] comp1540minVal;
    wire [5:0] comp1540minI, comp1540minJ;
    Comparator comp1540(SADValues[3172*12 +: 12], 49, 36, SADValues[3235*12 +: 12], 50, 35, comp1540minVal, comp1540minI, comp1540minJ);
    wire [11:0] comp1541minVal;
    wire [5:0] comp1541minI, comp1541minJ;
    Comparator comp1541(SADValues[3298*12 +: 12], 51, 34, SADValues[3361*12 +: 12], 52, 33, comp1541minVal, comp1541minI, comp1541minJ);
    wire [11:0] comp1542minVal;
    wire [5:0] comp1542minI, comp1542minJ;
    Comparator comp1542(SADValues[3424*12 +: 12], 53, 32, SADValues[3487*12 +: 12], 54, 31, comp1542minVal, comp1542minI, comp1542minJ);
    wire [11:0] comp1543minVal;
    wire [5:0] comp1543minI, comp1543minJ;
    Comparator comp1543(SADValues[3550*12 +: 12], 55, 30, SADValues[3613*12 +: 12], 56, 29, comp1543minVal, comp1543minI, comp1543minJ);
    wire [11:0] comp1544minVal;
    wire [5:0] comp1544minI, comp1544minJ;
    Comparator comp1544(SADValues[3676*12 +: 12], 57, 28, SADValues[3739*12 +: 12], 58, 27, comp1544minVal, comp1544minI, comp1544minJ);
    wire [11:0] comp1545minVal;
    wire [5:0] comp1545minI, comp1545minJ;
    Comparator comp1545(SADValues[3802*12 +: 12], 59, 26, SADValues[3865*12 +: 12], 60, 25, comp1545minVal, comp1545minI, comp1545minJ);
    wire [11:0] comp1546minVal;
    wire [5:0] comp1546minI, comp1546minJ;
    Comparator comp1546(SADValues[3866*12 +: 12], 60, 26, SADValues[3803*12 +: 12], 59, 27, comp1546minVal, comp1546minI, comp1546minJ);
    wire [11:0] comp1547minVal;
    wire [5:0] comp1547minI, comp1547minJ;
    Comparator comp1547(SADValues[3740*12 +: 12], 58, 28, SADValues[3677*12 +: 12], 57, 29, comp1547minVal, comp1547minI, comp1547minJ);
    wire [11:0] comp1548minVal;
    wire [5:0] comp1548minI, comp1548minJ;
    Comparator comp1548(SADValues[3614*12 +: 12], 56, 30, SADValues[3551*12 +: 12], 55, 31, comp1548minVal, comp1548minI, comp1548minJ);
    wire [11:0] comp1549minVal;
    wire [5:0] comp1549minI, comp1549minJ;
    Comparator comp1549(SADValues[3488*12 +: 12], 54, 32, SADValues[3425*12 +: 12], 53, 33, comp1549minVal, comp1549minI, comp1549minJ);
    wire [11:0] comp1550minVal;
    wire [5:0] comp1550minI, comp1550minJ;
    Comparator comp1550(SADValues[3362*12 +: 12], 52, 34, SADValues[3299*12 +: 12], 51, 35, comp1550minVal, comp1550minI, comp1550minJ);
    wire [11:0] comp1551minVal;
    wire [5:0] comp1551minI, comp1551minJ;
    Comparator comp1551(SADValues[3236*12 +: 12], 50, 36, SADValues[3173*12 +: 12], 49, 37, comp1551minVal, comp1551minI, comp1551minJ);
    wire [11:0] comp1552minVal;
    wire [5:0] comp1552minI, comp1552minJ;
    Comparator comp1552(SADValues[3110*12 +: 12], 48, 38, SADValues[3047*12 +: 12], 47, 39, comp1552minVal, comp1552minI, comp1552minJ);
    wire [11:0] comp1553minVal;
    wire [5:0] comp1553minI, comp1553minJ;
    Comparator comp1553(SADValues[2984*12 +: 12], 46, 40, SADValues[2921*12 +: 12], 45, 41, comp1553minVal, comp1553minI, comp1553minJ);
    wire [11:0] comp1554minVal;
    wire [5:0] comp1554minI, comp1554minJ;
    Comparator comp1554(SADValues[2858*12 +: 12], 44, 42, SADValues[2795*12 +: 12], 43, 43, comp1554minVal, comp1554minI, comp1554minJ);
    wire [11:0] comp1555minVal;
    wire [5:0] comp1555minI, comp1555minJ;
    Comparator comp1555(SADValues[2732*12 +: 12], 42, 44, SADValues[2669*12 +: 12], 41, 45, comp1555minVal, comp1555minI, comp1555minJ);
    wire [11:0] comp1556minVal;
    wire [5:0] comp1556minI, comp1556minJ;
    Comparator comp1556(SADValues[2606*12 +: 12], 40, 46, SADValues[2543*12 +: 12], 39, 47, comp1556minVal, comp1556minI, comp1556minJ);
    wire [11:0] comp1557minVal;
    wire [5:0] comp1557minI, comp1557minJ;
    Comparator comp1557(SADValues[2480*12 +: 12], 38, 48, SADValues[2417*12 +: 12], 37, 49, comp1557minVal, comp1557minI, comp1557minJ);
    wire [11:0] comp1558minVal;
    wire [5:0] comp1558minI, comp1558minJ;
    Comparator comp1558(SADValues[2354*12 +: 12], 36, 50, SADValues[2291*12 +: 12], 35, 51, comp1558minVal, comp1558minI, comp1558minJ);
    wire [11:0] comp1559minVal;
    wire [5:0] comp1559minI, comp1559minJ;
    Comparator comp1559(SADValues[2228*12 +: 12], 34, 52, SADValues[2165*12 +: 12], 33, 53, comp1559minVal, comp1559minI, comp1559minJ);
    wire [11:0] comp1560minVal;
    wire [5:0] comp1560minI, comp1560minJ;
    Comparator comp1560(SADValues[2102*12 +: 12], 32, 54, SADValues[2039*12 +: 12], 31, 55, comp1560minVal, comp1560minI, comp1560minJ);
    wire [11:0] comp1561minVal;
    wire [5:0] comp1561minI, comp1561minJ;
    Comparator comp1561(SADValues[1976*12 +: 12], 30, 56, SADValues[1913*12 +: 12], 29, 57, comp1561minVal, comp1561minI, comp1561minJ);
    wire [11:0] comp1562minVal;
    wire [5:0] comp1562minI, comp1562minJ;
    Comparator comp1562(SADValues[1850*12 +: 12], 28, 58, SADValues[1787*12 +: 12], 27, 59, comp1562minVal, comp1562minI, comp1562minJ);
    wire [11:0] comp1563minVal;
    wire [5:0] comp1563minI, comp1563minJ;
    Comparator comp1563(SADValues[1724*12 +: 12], 26, 60, SADValues[1788*12 +: 12], 27, 60, comp1563minVal, comp1563minI, comp1563minJ);
    wire [11:0] comp1564minVal;
    wire [5:0] comp1564minI, comp1564minJ;
    Comparator comp1564(SADValues[1851*12 +: 12], 28, 59, SADValues[1914*12 +: 12], 29, 58, comp1564minVal, comp1564minI, comp1564minJ);
    wire [11:0] comp1565minVal;
    wire [5:0] comp1565minI, comp1565minJ;
    Comparator comp1565(SADValues[1977*12 +: 12], 30, 57, SADValues[2040*12 +: 12], 31, 56, comp1565minVal, comp1565minI, comp1565minJ);
    wire [11:0] comp1566minVal;
    wire [5:0] comp1566minI, comp1566minJ;
    Comparator comp1566(SADValues[2103*12 +: 12], 32, 55, SADValues[2166*12 +: 12], 33, 54, comp1566minVal, comp1566minI, comp1566minJ);
    wire [11:0] comp1567minVal;
    wire [5:0] comp1567minI, comp1567minJ;
    Comparator comp1567(SADValues[2229*12 +: 12], 34, 53, SADValues[2292*12 +: 12], 35, 52, comp1567minVal, comp1567minI, comp1567minJ);
    wire [11:0] comp1568minVal;
    wire [5:0] comp1568minI, comp1568minJ;
    Comparator comp1568(SADValues[2355*12 +: 12], 36, 51, SADValues[2418*12 +: 12], 37, 50, comp1568minVal, comp1568minI, comp1568minJ);
    wire [11:0] comp1569minVal;
    wire [5:0] comp1569minI, comp1569minJ;
    Comparator comp1569(SADValues[2481*12 +: 12], 38, 49, SADValues[2544*12 +: 12], 39, 48, comp1569minVal, comp1569minI, comp1569minJ);
    wire [11:0] comp1570minVal;
    wire [5:0] comp1570minI, comp1570minJ;
    Comparator comp1570(SADValues[2607*12 +: 12], 40, 47, SADValues[2670*12 +: 12], 41, 46, comp1570minVal, comp1570minI, comp1570minJ);
    wire [11:0] comp1571minVal;
    wire [5:0] comp1571minI, comp1571minJ;
    Comparator comp1571(SADValues[2733*12 +: 12], 42, 45, SADValues[2796*12 +: 12], 43, 44, comp1571minVal, comp1571minI, comp1571minJ);
    wire [11:0] comp1572minVal;
    wire [5:0] comp1572minI, comp1572minJ;
    Comparator comp1572(SADValues[2859*12 +: 12], 44, 43, SADValues[2922*12 +: 12], 45, 42, comp1572minVal, comp1572minI, comp1572minJ);
    wire [11:0] comp1573minVal;
    wire [5:0] comp1573minI, comp1573minJ;
    Comparator comp1573(SADValues[2985*12 +: 12], 46, 41, SADValues[3048*12 +: 12], 47, 40, comp1573minVal, comp1573minI, comp1573minJ);
    wire [11:0] comp1574minVal;
    wire [5:0] comp1574minI, comp1574minJ;
    Comparator comp1574(SADValues[3111*12 +: 12], 48, 39, SADValues[3174*12 +: 12], 49, 38, comp1574minVal, comp1574minI, comp1574minJ);
    wire [11:0] comp1575minVal;
    wire [5:0] comp1575minI, comp1575minJ;
    Comparator comp1575(SADValues[3237*12 +: 12], 50, 37, SADValues[3300*12 +: 12], 51, 36, comp1575minVal, comp1575minI, comp1575minJ);
    wire [11:0] comp1576minVal;
    wire [5:0] comp1576minI, comp1576minJ;
    Comparator comp1576(SADValues[3363*12 +: 12], 52, 35, SADValues[3426*12 +: 12], 53, 34, comp1576minVal, comp1576minI, comp1576minJ);
    wire [11:0] comp1577minVal;
    wire [5:0] comp1577minI, comp1577minJ;
    Comparator comp1577(SADValues[3489*12 +: 12], 54, 33, SADValues[3552*12 +: 12], 55, 32, comp1577minVal, comp1577minI, comp1577minJ);
    wire [11:0] comp1578minVal;
    wire [5:0] comp1578minI, comp1578minJ;
    Comparator comp1578(SADValues[3615*12 +: 12], 56, 31, SADValues[3678*12 +: 12], 57, 30, comp1578minVal, comp1578minI, comp1578minJ);
    wire [11:0] comp1579minVal;
    wire [5:0] comp1579minI, comp1579minJ;
    Comparator comp1579(SADValues[3741*12 +: 12], 58, 29, SADValues[3804*12 +: 12], 59, 28, comp1579minVal, comp1579minI, comp1579minJ);
    wire [11:0] comp1580minVal;
    wire [5:0] comp1580minI, comp1580minJ;
    Comparator comp1580(SADValues[3867*12 +: 12], 60, 27, SADValues[3868*12 +: 12], 60, 28, comp1580minVal, comp1580minI, comp1580minJ);
    wire [11:0] comp1581minVal;
    wire [5:0] comp1581minI, comp1581minJ;
    Comparator comp1581(SADValues[3805*12 +: 12], 59, 29, SADValues[3742*12 +: 12], 58, 30, comp1581minVal, comp1581minI, comp1581minJ);
    wire [11:0] comp1582minVal;
    wire [5:0] comp1582minI, comp1582minJ;
    Comparator comp1582(SADValues[3679*12 +: 12], 57, 31, SADValues[3616*12 +: 12], 56, 32, comp1582minVal, comp1582minI, comp1582minJ);
    wire [11:0] comp1583minVal;
    wire [5:0] comp1583minI, comp1583minJ;
    Comparator comp1583(SADValues[3553*12 +: 12], 55, 33, SADValues[3490*12 +: 12], 54, 34, comp1583minVal, comp1583minI, comp1583minJ);
    wire [11:0] comp1584minVal;
    wire [5:0] comp1584minI, comp1584minJ;
    Comparator comp1584(SADValues[3427*12 +: 12], 53, 35, SADValues[3364*12 +: 12], 52, 36, comp1584minVal, comp1584minI, comp1584minJ);
    wire [11:0] comp1585minVal;
    wire [5:0] comp1585minI, comp1585minJ;
    Comparator comp1585(SADValues[3301*12 +: 12], 51, 37, SADValues[3238*12 +: 12], 50, 38, comp1585minVal, comp1585minI, comp1585minJ);
    wire [11:0] comp1586minVal;
    wire [5:0] comp1586minI, comp1586minJ;
    Comparator comp1586(SADValues[3175*12 +: 12], 49, 39, SADValues[3112*12 +: 12], 48, 40, comp1586minVal, comp1586minI, comp1586minJ);
    wire [11:0] comp1587minVal;
    wire [5:0] comp1587minI, comp1587minJ;
    Comparator comp1587(SADValues[3049*12 +: 12], 47, 41, SADValues[2986*12 +: 12], 46, 42, comp1587minVal, comp1587minI, comp1587minJ);
    wire [11:0] comp1588minVal;
    wire [5:0] comp1588minI, comp1588minJ;
    Comparator comp1588(SADValues[2923*12 +: 12], 45, 43, SADValues[2860*12 +: 12], 44, 44, comp1588minVal, comp1588minI, comp1588minJ);
    wire [11:0] comp1589minVal;
    wire [5:0] comp1589minI, comp1589minJ;
    Comparator comp1589(SADValues[2797*12 +: 12], 43, 45, SADValues[2734*12 +: 12], 42, 46, comp1589minVal, comp1589minI, comp1589minJ);
    wire [11:0] comp1590minVal;
    wire [5:0] comp1590minI, comp1590minJ;
    Comparator comp1590(SADValues[2671*12 +: 12], 41, 47, SADValues[2608*12 +: 12], 40, 48, comp1590minVal, comp1590minI, comp1590minJ);
    wire [11:0] comp1591minVal;
    wire [5:0] comp1591minI, comp1591minJ;
    Comparator comp1591(SADValues[2545*12 +: 12], 39, 49, SADValues[2482*12 +: 12], 38, 50, comp1591minVal, comp1591minI, comp1591minJ);
    wire [11:0] comp1592minVal;
    wire [5:0] comp1592minI, comp1592minJ;
    Comparator comp1592(SADValues[2419*12 +: 12], 37, 51, SADValues[2356*12 +: 12], 36, 52, comp1592minVal, comp1592minI, comp1592minJ);
    wire [11:0] comp1593minVal;
    wire [5:0] comp1593minI, comp1593minJ;
    Comparator comp1593(SADValues[2293*12 +: 12], 35, 53, SADValues[2230*12 +: 12], 34, 54, comp1593minVal, comp1593minI, comp1593minJ);
    wire [11:0] comp1594minVal;
    wire [5:0] comp1594minI, comp1594minJ;
    Comparator comp1594(SADValues[2167*12 +: 12], 33, 55, SADValues[2104*12 +: 12], 32, 56, comp1594minVal, comp1594minI, comp1594minJ);
    wire [11:0] comp1595minVal;
    wire [5:0] comp1595minI, comp1595minJ;
    Comparator comp1595(SADValues[2041*12 +: 12], 31, 57, SADValues[1978*12 +: 12], 30, 58, comp1595minVal, comp1595minI, comp1595minJ);
    wire [11:0] comp1596minVal;
    wire [5:0] comp1596minI, comp1596minJ;
    Comparator comp1596(SADValues[1915*12 +: 12], 29, 59, SADValues[1852*12 +: 12], 28, 60, comp1596minVal, comp1596minI, comp1596minJ);
    wire [11:0] comp1597minVal;
    wire [5:0] comp1597minI, comp1597minJ;
    Comparator comp1597(SADValues[1916*12 +: 12], 29, 60, SADValues[1979*12 +: 12], 30, 59, comp1597minVal, comp1597minI, comp1597minJ);
    wire [11:0] comp1598minVal;
    wire [5:0] comp1598minI, comp1598minJ;
    Comparator comp1598(SADValues[2042*12 +: 12], 31, 58, SADValues[2105*12 +: 12], 32, 57, comp1598minVal, comp1598minI, comp1598minJ);
    wire [11:0] comp1599minVal;
    wire [5:0] comp1599minI, comp1599minJ;
    Comparator comp1599(SADValues[2168*12 +: 12], 33, 56, SADValues[2231*12 +: 12], 34, 55, comp1599minVal, comp1599minI, comp1599minJ);
    wire [11:0] comp1600minVal;
    wire [5:0] comp1600minI, comp1600minJ;
    Comparator comp1600(SADValues[2294*12 +: 12], 35, 54, SADValues[2357*12 +: 12], 36, 53, comp1600minVal, comp1600minI, comp1600minJ);
    wire [11:0] comp1601minVal;
    wire [5:0] comp1601minI, comp1601minJ;
    Comparator comp1601(SADValues[2420*12 +: 12], 37, 52, SADValues[2483*12 +: 12], 38, 51, comp1601minVal, comp1601minI, comp1601minJ);
    wire [11:0] comp1602minVal;
    wire [5:0] comp1602minI, comp1602minJ;
    Comparator comp1602(SADValues[2546*12 +: 12], 39, 50, SADValues[2609*12 +: 12], 40, 49, comp1602minVal, comp1602minI, comp1602minJ);
    wire [11:0] comp1603minVal;
    wire [5:0] comp1603minI, comp1603minJ;
    Comparator comp1603(SADValues[2672*12 +: 12], 41, 48, SADValues[2735*12 +: 12], 42, 47, comp1603minVal, comp1603minI, comp1603minJ);
    wire [11:0] comp1604minVal;
    wire [5:0] comp1604minI, comp1604minJ;
    Comparator comp1604(SADValues[2798*12 +: 12], 43, 46, SADValues[2861*12 +: 12], 44, 45, comp1604minVal, comp1604minI, comp1604minJ);
    wire [11:0] comp1605minVal;
    wire [5:0] comp1605minI, comp1605minJ;
    Comparator comp1605(SADValues[2924*12 +: 12], 45, 44, SADValues[2987*12 +: 12], 46, 43, comp1605minVal, comp1605minI, comp1605minJ);
    wire [11:0] comp1606minVal;
    wire [5:0] comp1606minI, comp1606minJ;
    Comparator comp1606(SADValues[3050*12 +: 12], 47, 42, SADValues[3113*12 +: 12], 48, 41, comp1606minVal, comp1606minI, comp1606minJ);
    wire [11:0] comp1607minVal;
    wire [5:0] comp1607minI, comp1607minJ;
    Comparator comp1607(SADValues[3176*12 +: 12], 49, 40, SADValues[3239*12 +: 12], 50, 39, comp1607minVal, comp1607minI, comp1607minJ);
    wire [11:0] comp1608minVal;
    wire [5:0] comp1608minI, comp1608minJ;
    Comparator comp1608(SADValues[3302*12 +: 12], 51, 38, SADValues[3365*12 +: 12], 52, 37, comp1608minVal, comp1608minI, comp1608minJ);
    wire [11:0] comp1609minVal;
    wire [5:0] comp1609minI, comp1609minJ;
    Comparator comp1609(SADValues[3428*12 +: 12], 53, 36, SADValues[3491*12 +: 12], 54, 35, comp1609minVal, comp1609minI, comp1609minJ);
    wire [11:0] comp1610minVal;
    wire [5:0] comp1610minI, comp1610minJ;
    Comparator comp1610(SADValues[3554*12 +: 12], 55, 34, SADValues[3617*12 +: 12], 56, 33, comp1610minVal, comp1610minI, comp1610minJ);
    wire [11:0] comp1611minVal;
    wire [5:0] comp1611minI, comp1611minJ;
    Comparator comp1611(SADValues[3680*12 +: 12], 57, 32, SADValues[3743*12 +: 12], 58, 31, comp1611minVal, comp1611minI, comp1611minJ);
    wire [11:0] comp1612minVal;
    wire [5:0] comp1612minI, comp1612minJ;
    Comparator comp1612(SADValues[3806*12 +: 12], 59, 30, SADValues[3869*12 +: 12], 60, 29, comp1612minVal, comp1612minI, comp1612minJ);
    wire [11:0] comp1613minVal;
    wire [5:0] comp1613minI, comp1613minJ;
    Comparator comp1613(SADValues[3870*12 +: 12], 60, 30, SADValues[3807*12 +: 12], 59, 31, comp1613minVal, comp1613minI, comp1613minJ);
    wire [11:0] comp1614minVal;
    wire [5:0] comp1614minI, comp1614minJ;
    Comparator comp1614(SADValues[3744*12 +: 12], 58, 32, SADValues[3681*12 +: 12], 57, 33, comp1614minVal, comp1614minI, comp1614minJ);
    wire [11:0] comp1615minVal;
    wire [5:0] comp1615minI, comp1615minJ;
    Comparator comp1615(SADValues[3618*12 +: 12], 56, 34, SADValues[3555*12 +: 12], 55, 35, comp1615minVal, comp1615minI, comp1615minJ);
    wire [11:0] comp1616minVal;
    wire [5:0] comp1616minI, comp1616minJ;
    Comparator comp1616(SADValues[3492*12 +: 12], 54, 36, SADValues[3429*12 +: 12], 53, 37, comp1616minVal, comp1616minI, comp1616minJ);
    wire [11:0] comp1617minVal;
    wire [5:0] comp1617minI, comp1617minJ;
    Comparator comp1617(SADValues[3366*12 +: 12], 52, 38, SADValues[3303*12 +: 12], 51, 39, comp1617minVal, comp1617minI, comp1617minJ);
    wire [11:0] comp1618minVal;
    wire [5:0] comp1618minI, comp1618minJ;
    Comparator comp1618(SADValues[3240*12 +: 12], 50, 40, SADValues[3177*12 +: 12], 49, 41, comp1618minVal, comp1618minI, comp1618minJ);
    wire [11:0] comp1619minVal;
    wire [5:0] comp1619minI, comp1619minJ;
    Comparator comp1619(SADValues[3114*12 +: 12], 48, 42, SADValues[3051*12 +: 12], 47, 43, comp1619minVal, comp1619minI, comp1619minJ);
    wire [11:0] comp1620minVal;
    wire [5:0] comp1620minI, comp1620minJ;
    Comparator comp1620(SADValues[2988*12 +: 12], 46, 44, SADValues[2925*12 +: 12], 45, 45, comp1620minVal, comp1620minI, comp1620minJ);
    wire [11:0] comp1621minVal;
    wire [5:0] comp1621minI, comp1621minJ;
    Comparator comp1621(SADValues[2862*12 +: 12], 44, 46, SADValues[2799*12 +: 12], 43, 47, comp1621minVal, comp1621minI, comp1621minJ);
    wire [11:0] comp1622minVal;
    wire [5:0] comp1622minI, comp1622minJ;
    Comparator comp1622(SADValues[2736*12 +: 12], 42, 48, SADValues[2673*12 +: 12], 41, 49, comp1622minVal, comp1622minI, comp1622minJ);
    wire [11:0] comp1623minVal;
    wire [5:0] comp1623minI, comp1623minJ;
    Comparator comp1623(SADValues[2610*12 +: 12], 40, 50, SADValues[2547*12 +: 12], 39, 51, comp1623minVal, comp1623minI, comp1623minJ);
    wire [11:0] comp1624minVal;
    wire [5:0] comp1624minI, comp1624minJ;
    Comparator comp1624(SADValues[2484*12 +: 12], 38, 52, SADValues[2421*12 +: 12], 37, 53, comp1624minVal, comp1624minI, comp1624minJ);
    wire [11:0] comp1625minVal;
    wire [5:0] comp1625minI, comp1625minJ;
    Comparator comp1625(SADValues[2358*12 +: 12], 36, 54, SADValues[2295*12 +: 12], 35, 55, comp1625minVal, comp1625minI, comp1625minJ);
    wire [11:0] comp1626minVal;
    wire [5:0] comp1626minI, comp1626minJ;
    Comparator comp1626(SADValues[2232*12 +: 12], 34, 56, SADValues[2169*12 +: 12], 33, 57, comp1626minVal, comp1626minI, comp1626minJ);
    wire [11:0] comp1627minVal;
    wire [5:0] comp1627minI, comp1627minJ;
    Comparator comp1627(SADValues[2106*12 +: 12], 32, 58, SADValues[2043*12 +: 12], 31, 59, comp1627minVal, comp1627minI, comp1627minJ);
    wire [11:0] comp1628minVal;
    wire [5:0] comp1628minI, comp1628minJ;
    Comparator comp1628(SADValues[1980*12 +: 12], 30, 60, SADValues[2044*12 +: 12], 31, 60, comp1628minVal, comp1628minI, comp1628minJ);
    wire [11:0] comp1629minVal;
    wire [5:0] comp1629minI, comp1629minJ;
    Comparator comp1629(SADValues[2107*12 +: 12], 32, 59, SADValues[2170*12 +: 12], 33, 58, comp1629minVal, comp1629minI, comp1629minJ);
    wire [11:0] comp1630minVal;
    wire [5:0] comp1630minI, comp1630minJ;
    Comparator comp1630(SADValues[2233*12 +: 12], 34, 57, SADValues[2296*12 +: 12], 35, 56, comp1630minVal, comp1630minI, comp1630minJ);
    wire [11:0] comp1631minVal;
    wire [5:0] comp1631minI, comp1631minJ;
    Comparator comp1631(SADValues[2359*12 +: 12], 36, 55, SADValues[2422*12 +: 12], 37, 54, comp1631minVal, comp1631minI, comp1631minJ);
    wire [11:0] comp1632minVal;
    wire [5:0] comp1632minI, comp1632minJ;
    Comparator comp1632(SADValues[2485*12 +: 12], 38, 53, SADValues[2548*12 +: 12], 39, 52, comp1632minVal, comp1632minI, comp1632minJ);
    wire [11:0] comp1633minVal;
    wire [5:0] comp1633minI, comp1633minJ;
    Comparator comp1633(SADValues[2611*12 +: 12], 40, 51, SADValues[2674*12 +: 12], 41, 50, comp1633minVal, comp1633minI, comp1633minJ);
    wire [11:0] comp1634minVal;
    wire [5:0] comp1634minI, comp1634minJ;
    Comparator comp1634(SADValues[2737*12 +: 12], 42, 49, SADValues[2800*12 +: 12], 43, 48, comp1634minVal, comp1634minI, comp1634minJ);
    wire [11:0] comp1635minVal;
    wire [5:0] comp1635minI, comp1635minJ;
    Comparator comp1635(SADValues[2863*12 +: 12], 44, 47, SADValues[2926*12 +: 12], 45, 46, comp1635minVal, comp1635minI, comp1635minJ);
    wire [11:0] comp1636minVal;
    wire [5:0] comp1636minI, comp1636minJ;
    Comparator comp1636(SADValues[2989*12 +: 12], 46, 45, SADValues[3052*12 +: 12], 47, 44, comp1636minVal, comp1636minI, comp1636minJ);
    wire [11:0] comp1637minVal;
    wire [5:0] comp1637minI, comp1637minJ;
    Comparator comp1637(SADValues[3115*12 +: 12], 48, 43, SADValues[3178*12 +: 12], 49, 42, comp1637minVal, comp1637minI, comp1637minJ);
    wire [11:0] comp1638minVal;
    wire [5:0] comp1638minI, comp1638minJ;
    Comparator comp1638(SADValues[3241*12 +: 12], 50, 41, SADValues[3304*12 +: 12], 51, 40, comp1638minVal, comp1638minI, comp1638minJ);
    wire [11:0] comp1639minVal;
    wire [5:0] comp1639minI, comp1639minJ;
    Comparator comp1639(SADValues[3367*12 +: 12], 52, 39, SADValues[3430*12 +: 12], 53, 38, comp1639minVal, comp1639minI, comp1639minJ);
    wire [11:0] comp1640minVal;
    wire [5:0] comp1640minI, comp1640minJ;
    Comparator comp1640(SADValues[3493*12 +: 12], 54, 37, SADValues[3556*12 +: 12], 55, 36, comp1640minVal, comp1640minI, comp1640minJ);
    wire [11:0] comp1641minVal;
    wire [5:0] comp1641minI, comp1641minJ;
    Comparator comp1641(SADValues[3619*12 +: 12], 56, 35, SADValues[3682*12 +: 12], 57, 34, comp1641minVal, comp1641minI, comp1641minJ);
    wire [11:0] comp1642minVal;
    wire [5:0] comp1642minI, comp1642minJ;
    Comparator comp1642(SADValues[3745*12 +: 12], 58, 33, SADValues[3808*12 +: 12], 59, 32, comp1642minVal, comp1642minI, comp1642minJ);
    wire [11:0] comp1643minVal;
    wire [5:0] comp1643minI, comp1643minJ;
    Comparator comp1643(SADValues[3871*12 +: 12], 60, 31, SADValues[3872*12 +: 12], 60, 32, comp1643minVal, comp1643minI, comp1643minJ);
    wire [11:0] comp1644minVal;
    wire [5:0] comp1644minI, comp1644minJ;
    Comparator comp1644(SADValues[3809*12 +: 12], 59, 33, SADValues[3746*12 +: 12], 58, 34, comp1644minVal, comp1644minI, comp1644minJ);
    wire [11:0] comp1645minVal;
    wire [5:0] comp1645minI, comp1645minJ;
    Comparator comp1645(SADValues[3683*12 +: 12], 57, 35, SADValues[3620*12 +: 12], 56, 36, comp1645minVal, comp1645minI, comp1645minJ);
    wire [11:0] comp1646minVal;
    wire [5:0] comp1646minI, comp1646minJ;
    Comparator comp1646(SADValues[3557*12 +: 12], 55, 37, SADValues[3494*12 +: 12], 54, 38, comp1646minVal, comp1646minI, comp1646minJ);
    wire [11:0] comp1647minVal;
    wire [5:0] comp1647minI, comp1647minJ;
    Comparator comp1647(SADValues[3431*12 +: 12], 53, 39, SADValues[3368*12 +: 12], 52, 40, comp1647minVal, comp1647minI, comp1647minJ);
    wire [11:0] comp1648minVal;
    wire [5:0] comp1648minI, comp1648minJ;
    Comparator comp1648(SADValues[3305*12 +: 12], 51, 41, SADValues[3242*12 +: 12], 50, 42, comp1648minVal, comp1648minI, comp1648minJ);
    wire [11:0] comp1649minVal;
    wire [5:0] comp1649minI, comp1649minJ;
    Comparator comp1649(SADValues[3179*12 +: 12], 49, 43, SADValues[3116*12 +: 12], 48, 44, comp1649minVal, comp1649minI, comp1649minJ);
    wire [11:0] comp1650minVal;
    wire [5:0] comp1650minI, comp1650minJ;
    Comparator comp1650(SADValues[3053*12 +: 12], 47, 45, SADValues[2990*12 +: 12], 46, 46, comp1650minVal, comp1650minI, comp1650minJ);
    wire [11:0] comp1651minVal;
    wire [5:0] comp1651minI, comp1651minJ;
    Comparator comp1651(SADValues[2927*12 +: 12], 45, 47, SADValues[2864*12 +: 12], 44, 48, comp1651minVal, comp1651minI, comp1651minJ);
    wire [11:0] comp1652minVal;
    wire [5:0] comp1652minI, comp1652minJ;
    Comparator comp1652(SADValues[2801*12 +: 12], 43, 49, SADValues[2738*12 +: 12], 42, 50, comp1652minVal, comp1652minI, comp1652minJ);
    wire [11:0] comp1653minVal;
    wire [5:0] comp1653minI, comp1653minJ;
    Comparator comp1653(SADValues[2675*12 +: 12], 41, 51, SADValues[2612*12 +: 12], 40, 52, comp1653minVal, comp1653minI, comp1653minJ);
    wire [11:0] comp1654minVal;
    wire [5:0] comp1654minI, comp1654minJ;
    Comparator comp1654(SADValues[2549*12 +: 12], 39, 53, SADValues[2486*12 +: 12], 38, 54, comp1654minVal, comp1654minI, comp1654minJ);
    wire [11:0] comp1655minVal;
    wire [5:0] comp1655minI, comp1655minJ;
    Comparator comp1655(SADValues[2423*12 +: 12], 37, 55, SADValues[2360*12 +: 12], 36, 56, comp1655minVal, comp1655minI, comp1655minJ);
    wire [11:0] comp1656minVal;
    wire [5:0] comp1656minI, comp1656minJ;
    Comparator comp1656(SADValues[2297*12 +: 12], 35, 57, SADValues[2234*12 +: 12], 34, 58, comp1656minVal, comp1656minI, comp1656minJ);
    wire [11:0] comp1657minVal;
    wire [5:0] comp1657minI, comp1657minJ;
    Comparator comp1657(SADValues[2171*12 +: 12], 33, 59, SADValues[2108*12 +: 12], 32, 60, comp1657minVal, comp1657minI, comp1657minJ);
    wire [11:0] comp1658minVal;
    wire [5:0] comp1658minI, comp1658minJ;
    Comparator comp1658(SADValues[2172*12 +: 12], 33, 60, SADValues[2235*12 +: 12], 34, 59, comp1658minVal, comp1658minI, comp1658minJ);
    wire [11:0] comp1659minVal;
    wire [5:0] comp1659minI, comp1659minJ;
    Comparator comp1659(SADValues[2298*12 +: 12], 35, 58, SADValues[2361*12 +: 12], 36, 57, comp1659minVal, comp1659minI, comp1659minJ);
    wire [11:0] comp1660minVal;
    wire [5:0] comp1660minI, comp1660minJ;
    Comparator comp1660(SADValues[2424*12 +: 12], 37, 56, SADValues[2487*12 +: 12], 38, 55, comp1660minVal, comp1660minI, comp1660minJ);
    wire [11:0] comp1661minVal;
    wire [5:0] comp1661minI, comp1661minJ;
    Comparator comp1661(SADValues[2550*12 +: 12], 39, 54, SADValues[2613*12 +: 12], 40, 53, comp1661minVal, comp1661minI, comp1661minJ);
    wire [11:0] comp1662minVal;
    wire [5:0] comp1662minI, comp1662minJ;
    Comparator comp1662(SADValues[2676*12 +: 12], 41, 52, SADValues[2739*12 +: 12], 42, 51, comp1662minVal, comp1662minI, comp1662minJ);
    wire [11:0] comp1663minVal;
    wire [5:0] comp1663minI, comp1663minJ;
    Comparator comp1663(SADValues[2802*12 +: 12], 43, 50, SADValues[2865*12 +: 12], 44, 49, comp1663minVal, comp1663minI, comp1663minJ);
    wire [11:0] comp1664minVal;
    wire [5:0] comp1664minI, comp1664minJ;
    Comparator comp1664(SADValues[2928*12 +: 12], 45, 48, SADValues[2991*12 +: 12], 46, 47, comp1664minVal, comp1664minI, comp1664minJ);
    wire [11:0] comp1665minVal;
    wire [5:0] comp1665minI, comp1665minJ;
    Comparator comp1665(SADValues[3054*12 +: 12], 47, 46, SADValues[3117*12 +: 12], 48, 45, comp1665minVal, comp1665minI, comp1665minJ);
    wire [11:0] comp1666minVal;
    wire [5:0] comp1666minI, comp1666minJ;
    Comparator comp1666(SADValues[3180*12 +: 12], 49, 44, SADValues[3243*12 +: 12], 50, 43, comp1666minVal, comp1666minI, comp1666minJ);
    wire [11:0] comp1667minVal;
    wire [5:0] comp1667minI, comp1667minJ;
    Comparator comp1667(SADValues[3306*12 +: 12], 51, 42, SADValues[3369*12 +: 12], 52, 41, comp1667minVal, comp1667minI, comp1667minJ);
    wire [11:0] comp1668minVal;
    wire [5:0] comp1668minI, comp1668minJ;
    Comparator comp1668(SADValues[3432*12 +: 12], 53, 40, SADValues[3495*12 +: 12], 54, 39, comp1668minVal, comp1668minI, comp1668minJ);
    wire [11:0] comp1669minVal;
    wire [5:0] comp1669minI, comp1669minJ;
    Comparator comp1669(SADValues[3558*12 +: 12], 55, 38, SADValues[3621*12 +: 12], 56, 37, comp1669minVal, comp1669minI, comp1669minJ);
    wire [11:0] comp1670minVal;
    wire [5:0] comp1670minI, comp1670minJ;
    Comparator comp1670(SADValues[3684*12 +: 12], 57, 36, SADValues[3747*12 +: 12], 58, 35, comp1670minVal, comp1670minI, comp1670minJ);
    wire [11:0] comp1671minVal;
    wire [5:0] comp1671minI, comp1671minJ;
    Comparator comp1671(SADValues[3810*12 +: 12], 59, 34, SADValues[3873*12 +: 12], 60, 33, comp1671minVal, comp1671minI, comp1671minJ);
    wire [11:0] comp1672minVal;
    wire [5:0] comp1672minI, comp1672minJ;
    Comparator comp1672(SADValues[3874*12 +: 12], 60, 34, SADValues[3811*12 +: 12], 59, 35, comp1672minVal, comp1672minI, comp1672minJ);
    wire [11:0] comp1673minVal;
    wire [5:0] comp1673minI, comp1673minJ;
    Comparator comp1673(SADValues[3748*12 +: 12], 58, 36, SADValues[3685*12 +: 12], 57, 37, comp1673minVal, comp1673minI, comp1673minJ);
    wire [11:0] comp1674minVal;
    wire [5:0] comp1674minI, comp1674minJ;
    Comparator comp1674(SADValues[3622*12 +: 12], 56, 38, SADValues[3559*12 +: 12], 55, 39, comp1674minVal, comp1674minI, comp1674minJ);
    wire [11:0] comp1675minVal;
    wire [5:0] comp1675minI, comp1675minJ;
    Comparator comp1675(SADValues[3496*12 +: 12], 54, 40, SADValues[3433*12 +: 12], 53, 41, comp1675minVal, comp1675minI, comp1675minJ);
    wire [11:0] comp1676minVal;
    wire [5:0] comp1676minI, comp1676minJ;
    Comparator comp1676(SADValues[3370*12 +: 12], 52, 42, SADValues[3307*12 +: 12], 51, 43, comp1676minVal, comp1676minI, comp1676minJ);
    wire [11:0] comp1677minVal;
    wire [5:0] comp1677minI, comp1677minJ;
    Comparator comp1677(SADValues[3244*12 +: 12], 50, 44, SADValues[3181*12 +: 12], 49, 45, comp1677minVal, comp1677minI, comp1677minJ);
    wire [11:0] comp1678minVal;
    wire [5:0] comp1678minI, comp1678minJ;
    Comparator comp1678(SADValues[3118*12 +: 12], 48, 46, SADValues[3055*12 +: 12], 47, 47, comp1678minVal, comp1678minI, comp1678minJ);
    wire [11:0] comp1679minVal;
    wire [5:0] comp1679minI, comp1679minJ;
    Comparator comp1679(SADValues[2992*12 +: 12], 46, 48, SADValues[2929*12 +: 12], 45, 49, comp1679minVal, comp1679minI, comp1679minJ);
    wire [11:0] comp1680minVal;
    wire [5:0] comp1680minI, comp1680minJ;
    Comparator comp1680(SADValues[2866*12 +: 12], 44, 50, SADValues[2803*12 +: 12], 43, 51, comp1680minVal, comp1680minI, comp1680minJ);
    wire [11:0] comp1681minVal;
    wire [5:0] comp1681minI, comp1681minJ;
    Comparator comp1681(SADValues[2740*12 +: 12], 42, 52, SADValues[2677*12 +: 12], 41, 53, comp1681minVal, comp1681minI, comp1681minJ);
    wire [11:0] comp1682minVal;
    wire [5:0] comp1682minI, comp1682minJ;
    Comparator comp1682(SADValues[2614*12 +: 12], 40, 54, SADValues[2551*12 +: 12], 39, 55, comp1682minVal, comp1682minI, comp1682minJ);
    wire [11:0] comp1683minVal;
    wire [5:0] comp1683minI, comp1683minJ;
    Comparator comp1683(SADValues[2488*12 +: 12], 38, 56, SADValues[2425*12 +: 12], 37, 57, comp1683minVal, comp1683minI, comp1683minJ);
    wire [11:0] comp1684minVal;
    wire [5:0] comp1684minI, comp1684minJ;
    Comparator comp1684(SADValues[2362*12 +: 12], 36, 58, SADValues[2299*12 +: 12], 35, 59, comp1684minVal, comp1684minI, comp1684minJ);
    wire [11:0] comp1685minVal;
    wire [5:0] comp1685minI, comp1685minJ;
    Comparator comp1685(SADValues[2236*12 +: 12], 34, 60, SADValues[2300*12 +: 12], 35, 60, comp1685minVal, comp1685minI, comp1685minJ);
    wire [11:0] comp1686minVal;
    wire [5:0] comp1686minI, comp1686minJ;
    Comparator comp1686(SADValues[2363*12 +: 12], 36, 59, SADValues[2426*12 +: 12], 37, 58, comp1686minVal, comp1686minI, comp1686minJ);
    wire [11:0] comp1687minVal;
    wire [5:0] comp1687minI, comp1687minJ;
    Comparator comp1687(SADValues[2489*12 +: 12], 38, 57, SADValues[2552*12 +: 12], 39, 56, comp1687minVal, comp1687minI, comp1687minJ);
    wire [11:0] comp1688minVal;
    wire [5:0] comp1688minI, comp1688minJ;
    Comparator comp1688(SADValues[2615*12 +: 12], 40, 55, SADValues[2678*12 +: 12], 41, 54, comp1688minVal, comp1688minI, comp1688minJ);
    wire [11:0] comp1689minVal;
    wire [5:0] comp1689minI, comp1689minJ;
    Comparator comp1689(SADValues[2741*12 +: 12], 42, 53, SADValues[2804*12 +: 12], 43, 52, comp1689minVal, comp1689minI, comp1689minJ);
    wire [11:0] comp1690minVal;
    wire [5:0] comp1690minI, comp1690minJ;
    Comparator comp1690(SADValues[2867*12 +: 12], 44, 51, SADValues[2930*12 +: 12], 45, 50, comp1690minVal, comp1690minI, comp1690minJ);
    wire [11:0] comp1691minVal;
    wire [5:0] comp1691minI, comp1691minJ;
    Comparator comp1691(SADValues[2993*12 +: 12], 46, 49, SADValues[3056*12 +: 12], 47, 48, comp1691minVal, comp1691minI, comp1691minJ);
    wire [11:0] comp1692minVal;
    wire [5:0] comp1692minI, comp1692minJ;
    Comparator comp1692(SADValues[3119*12 +: 12], 48, 47, SADValues[3182*12 +: 12], 49, 46, comp1692minVal, comp1692minI, comp1692minJ);
    wire [11:0] comp1693minVal;
    wire [5:0] comp1693minI, comp1693minJ;
    Comparator comp1693(SADValues[3245*12 +: 12], 50, 45, SADValues[3308*12 +: 12], 51, 44, comp1693minVal, comp1693minI, comp1693minJ);
    wire [11:0] comp1694minVal;
    wire [5:0] comp1694minI, comp1694minJ;
    Comparator comp1694(SADValues[3371*12 +: 12], 52, 43, SADValues[3434*12 +: 12], 53, 42, comp1694minVal, comp1694minI, comp1694minJ);
    wire [11:0] comp1695minVal;
    wire [5:0] comp1695minI, comp1695minJ;
    Comparator comp1695(SADValues[3497*12 +: 12], 54, 41, SADValues[3560*12 +: 12], 55, 40, comp1695minVal, comp1695minI, comp1695minJ);
    wire [11:0] comp1696minVal;
    wire [5:0] comp1696minI, comp1696minJ;
    Comparator comp1696(SADValues[3623*12 +: 12], 56, 39, SADValues[3686*12 +: 12], 57, 38, comp1696minVal, comp1696minI, comp1696minJ);
    wire [11:0] comp1697minVal;
    wire [5:0] comp1697minI, comp1697minJ;
    Comparator comp1697(SADValues[3749*12 +: 12], 58, 37, SADValues[3812*12 +: 12], 59, 36, comp1697minVal, comp1697minI, comp1697minJ);
    wire [11:0] comp1698minVal;
    wire [5:0] comp1698minI, comp1698minJ;
    Comparator comp1698(SADValues[3875*12 +: 12], 60, 35, SADValues[3876*12 +: 12], 60, 36, comp1698minVal, comp1698minI, comp1698minJ);
    wire [11:0] comp1699minVal;
    wire [5:0] comp1699minI, comp1699minJ;
    Comparator comp1699(SADValues[3813*12 +: 12], 59, 37, SADValues[3750*12 +: 12], 58, 38, comp1699minVal, comp1699minI, comp1699minJ);
    wire [11:0] comp1700minVal;
    wire [5:0] comp1700minI, comp1700minJ;
    Comparator comp1700(SADValues[3687*12 +: 12], 57, 39, SADValues[3624*12 +: 12], 56, 40, comp1700minVal, comp1700minI, comp1700minJ);
    wire [11:0] comp1701minVal;
    wire [5:0] comp1701minI, comp1701minJ;
    Comparator comp1701(SADValues[3561*12 +: 12], 55, 41, SADValues[3498*12 +: 12], 54, 42, comp1701minVal, comp1701minI, comp1701minJ);
    wire [11:0] comp1702minVal;
    wire [5:0] comp1702minI, comp1702minJ;
    Comparator comp1702(SADValues[3435*12 +: 12], 53, 43, SADValues[3372*12 +: 12], 52, 44, comp1702minVal, comp1702minI, comp1702minJ);
    wire [11:0] comp1703minVal;
    wire [5:0] comp1703minI, comp1703minJ;
    Comparator comp1703(SADValues[3309*12 +: 12], 51, 45, SADValues[3246*12 +: 12], 50, 46, comp1703minVal, comp1703minI, comp1703minJ);
    wire [11:0] comp1704minVal;
    wire [5:0] comp1704minI, comp1704minJ;
    Comparator comp1704(SADValues[3183*12 +: 12], 49, 47, SADValues[3120*12 +: 12], 48, 48, comp1704minVal, comp1704minI, comp1704minJ);
    wire [11:0] comp1705minVal;
    wire [5:0] comp1705minI, comp1705minJ;
    Comparator comp1705(SADValues[3057*12 +: 12], 47, 49, SADValues[2994*12 +: 12], 46, 50, comp1705minVal, comp1705minI, comp1705minJ);
    wire [11:0] comp1706minVal;
    wire [5:0] comp1706minI, comp1706minJ;
    Comparator comp1706(SADValues[2931*12 +: 12], 45, 51, SADValues[2868*12 +: 12], 44, 52, comp1706minVal, comp1706minI, comp1706minJ);
    wire [11:0] comp1707minVal;
    wire [5:0] comp1707minI, comp1707minJ;
    Comparator comp1707(SADValues[2805*12 +: 12], 43, 53, SADValues[2742*12 +: 12], 42, 54, comp1707minVal, comp1707minI, comp1707minJ);
    wire [11:0] comp1708minVal;
    wire [5:0] comp1708minI, comp1708minJ;
    Comparator comp1708(SADValues[2679*12 +: 12], 41, 55, SADValues[2616*12 +: 12], 40, 56, comp1708minVal, comp1708minI, comp1708minJ);
    wire [11:0] comp1709minVal;
    wire [5:0] comp1709minI, comp1709minJ;
    Comparator comp1709(SADValues[2553*12 +: 12], 39, 57, SADValues[2490*12 +: 12], 38, 58, comp1709minVal, comp1709minI, comp1709minJ);
    wire [11:0] comp1710minVal;
    wire [5:0] comp1710minI, comp1710minJ;
    Comparator comp1710(SADValues[2427*12 +: 12], 37, 59, SADValues[2364*12 +: 12], 36, 60, comp1710minVal, comp1710minI, comp1710minJ);
    wire [11:0] comp1711minVal;
    wire [5:0] comp1711minI, comp1711minJ;
    Comparator comp1711(SADValues[2428*12 +: 12], 37, 60, SADValues[2491*12 +: 12], 38, 59, comp1711minVal, comp1711minI, comp1711minJ);
    wire [11:0] comp1712minVal;
    wire [5:0] comp1712minI, comp1712minJ;
    Comparator comp1712(SADValues[2554*12 +: 12], 39, 58, SADValues[2617*12 +: 12], 40, 57, comp1712minVal, comp1712minI, comp1712minJ);
    wire [11:0] comp1713minVal;
    wire [5:0] comp1713minI, comp1713minJ;
    Comparator comp1713(SADValues[2680*12 +: 12], 41, 56, SADValues[2743*12 +: 12], 42, 55, comp1713minVal, comp1713minI, comp1713minJ);
    wire [11:0] comp1714minVal;
    wire [5:0] comp1714minI, comp1714minJ;
    Comparator comp1714(SADValues[2806*12 +: 12], 43, 54, SADValues[2869*12 +: 12], 44, 53, comp1714minVal, comp1714minI, comp1714minJ);
    wire [11:0] comp1715minVal;
    wire [5:0] comp1715minI, comp1715minJ;
    Comparator comp1715(SADValues[2932*12 +: 12], 45, 52, SADValues[2995*12 +: 12], 46, 51, comp1715minVal, comp1715minI, comp1715minJ);
    wire [11:0] comp1716minVal;
    wire [5:0] comp1716minI, comp1716minJ;
    Comparator comp1716(SADValues[3058*12 +: 12], 47, 50, SADValues[3121*12 +: 12], 48, 49, comp1716minVal, comp1716minI, comp1716minJ);
    wire [11:0] comp1717minVal;
    wire [5:0] comp1717minI, comp1717minJ;
    Comparator comp1717(SADValues[3184*12 +: 12], 49, 48, SADValues[3247*12 +: 12], 50, 47, comp1717minVal, comp1717minI, comp1717minJ);
    wire [11:0] comp1718minVal;
    wire [5:0] comp1718minI, comp1718minJ;
    Comparator comp1718(SADValues[3310*12 +: 12], 51, 46, SADValues[3373*12 +: 12], 52, 45, comp1718minVal, comp1718minI, comp1718minJ);
    wire [11:0] comp1719minVal;
    wire [5:0] comp1719minI, comp1719minJ;
    Comparator comp1719(SADValues[3436*12 +: 12], 53, 44, SADValues[3499*12 +: 12], 54, 43, comp1719minVal, comp1719minI, comp1719minJ);
    wire [11:0] comp1720minVal;
    wire [5:0] comp1720minI, comp1720minJ;
    Comparator comp1720(SADValues[3562*12 +: 12], 55, 42, SADValues[3625*12 +: 12], 56, 41, comp1720minVal, comp1720minI, comp1720minJ);
    wire [11:0] comp1721minVal;
    wire [5:0] comp1721minI, comp1721minJ;
    Comparator comp1721(SADValues[3688*12 +: 12], 57, 40, SADValues[3751*12 +: 12], 58, 39, comp1721minVal, comp1721minI, comp1721minJ);
    wire [11:0] comp1722minVal;
    wire [5:0] comp1722minI, comp1722minJ;
    Comparator comp1722(SADValues[3814*12 +: 12], 59, 38, SADValues[3877*12 +: 12], 60, 37, comp1722minVal, comp1722minI, comp1722minJ);
    wire [11:0] comp1723minVal;
    wire [5:0] comp1723minI, comp1723minJ;
    Comparator comp1723(SADValues[3878*12 +: 12], 60, 38, SADValues[3815*12 +: 12], 59, 39, comp1723minVal, comp1723minI, comp1723minJ);
    wire [11:0] comp1724minVal;
    wire [5:0] comp1724minI, comp1724minJ;
    Comparator comp1724(SADValues[3752*12 +: 12], 58, 40, SADValues[3689*12 +: 12], 57, 41, comp1724minVal, comp1724minI, comp1724minJ);
    wire [11:0] comp1725minVal;
    wire [5:0] comp1725minI, comp1725minJ;
    Comparator comp1725(SADValues[3626*12 +: 12], 56, 42, SADValues[3563*12 +: 12], 55, 43, comp1725minVal, comp1725minI, comp1725minJ);
    wire [11:0] comp1726minVal;
    wire [5:0] comp1726minI, comp1726minJ;
    Comparator comp1726(SADValues[3500*12 +: 12], 54, 44, SADValues[3437*12 +: 12], 53, 45, comp1726minVal, comp1726minI, comp1726minJ);
    wire [11:0] comp1727minVal;
    wire [5:0] comp1727minI, comp1727minJ;
    Comparator comp1727(SADValues[3374*12 +: 12], 52, 46, SADValues[3311*12 +: 12], 51, 47, comp1727minVal, comp1727minI, comp1727minJ);
    wire [11:0] comp1728minVal;
    wire [5:0] comp1728minI, comp1728minJ;
    Comparator comp1728(SADValues[3248*12 +: 12], 50, 48, SADValues[3185*12 +: 12], 49, 49, comp1728minVal, comp1728minI, comp1728minJ);
    wire [11:0] comp1729minVal;
    wire [5:0] comp1729minI, comp1729minJ;
    Comparator comp1729(SADValues[3122*12 +: 12], 48, 50, SADValues[3059*12 +: 12], 47, 51, comp1729minVal, comp1729minI, comp1729minJ);
    wire [11:0] comp1730minVal;
    wire [5:0] comp1730minI, comp1730minJ;
    Comparator comp1730(SADValues[2996*12 +: 12], 46, 52, SADValues[2933*12 +: 12], 45, 53, comp1730minVal, comp1730minI, comp1730minJ);
    wire [11:0] comp1731minVal;
    wire [5:0] comp1731minI, comp1731minJ;
    Comparator comp1731(SADValues[2870*12 +: 12], 44, 54, SADValues[2807*12 +: 12], 43, 55, comp1731minVal, comp1731minI, comp1731minJ);
    wire [11:0] comp1732minVal;
    wire [5:0] comp1732minI, comp1732minJ;
    Comparator comp1732(SADValues[2744*12 +: 12], 42, 56, SADValues[2681*12 +: 12], 41, 57, comp1732minVal, comp1732minI, comp1732minJ);
    wire [11:0] comp1733minVal;
    wire [5:0] comp1733minI, comp1733minJ;
    Comparator comp1733(SADValues[2618*12 +: 12], 40, 58, SADValues[2555*12 +: 12], 39, 59, comp1733minVal, comp1733minI, comp1733minJ);
    wire [11:0] comp1734minVal;
    wire [5:0] comp1734minI, comp1734minJ;
    Comparator comp1734(SADValues[2492*12 +: 12], 38, 60, SADValues[2556*12 +: 12], 39, 60, comp1734minVal, comp1734minI, comp1734minJ);
    wire [11:0] comp1735minVal;
    wire [5:0] comp1735minI, comp1735minJ;
    Comparator comp1735(SADValues[2619*12 +: 12], 40, 59, SADValues[2682*12 +: 12], 41, 58, comp1735minVal, comp1735minI, comp1735minJ);
    wire [11:0] comp1736minVal;
    wire [5:0] comp1736minI, comp1736minJ;
    Comparator comp1736(SADValues[2745*12 +: 12], 42, 57, SADValues[2808*12 +: 12], 43, 56, comp1736minVal, comp1736minI, comp1736minJ);
    wire [11:0] comp1737minVal;
    wire [5:0] comp1737minI, comp1737minJ;
    Comparator comp1737(SADValues[2871*12 +: 12], 44, 55, SADValues[2934*12 +: 12], 45, 54, comp1737minVal, comp1737minI, comp1737minJ);
    wire [11:0] comp1738minVal;
    wire [5:0] comp1738minI, comp1738minJ;
    Comparator comp1738(SADValues[2997*12 +: 12], 46, 53, SADValues[3060*12 +: 12], 47, 52, comp1738minVal, comp1738minI, comp1738minJ);
    wire [11:0] comp1739minVal;
    wire [5:0] comp1739minI, comp1739minJ;
    Comparator comp1739(SADValues[3123*12 +: 12], 48, 51, SADValues[3186*12 +: 12], 49, 50, comp1739minVal, comp1739minI, comp1739minJ);
    wire [11:0] comp1740minVal;
    wire [5:0] comp1740minI, comp1740minJ;
    Comparator comp1740(SADValues[3249*12 +: 12], 50, 49, SADValues[3312*12 +: 12], 51, 48, comp1740minVal, comp1740minI, comp1740minJ);
    wire [11:0] comp1741minVal;
    wire [5:0] comp1741minI, comp1741minJ;
    Comparator comp1741(SADValues[3375*12 +: 12], 52, 47, SADValues[3438*12 +: 12], 53, 46, comp1741minVal, comp1741minI, comp1741minJ);
    wire [11:0] comp1742minVal;
    wire [5:0] comp1742minI, comp1742minJ;
    Comparator comp1742(SADValues[3501*12 +: 12], 54, 45, SADValues[3564*12 +: 12], 55, 44, comp1742minVal, comp1742minI, comp1742minJ);
    wire [11:0] comp1743minVal;
    wire [5:0] comp1743minI, comp1743minJ;
    Comparator comp1743(SADValues[3627*12 +: 12], 56, 43, SADValues[3690*12 +: 12], 57, 42, comp1743minVal, comp1743minI, comp1743minJ);
    wire [11:0] comp1744minVal;
    wire [5:0] comp1744minI, comp1744minJ;
    Comparator comp1744(SADValues[3753*12 +: 12], 58, 41, SADValues[3816*12 +: 12], 59, 40, comp1744minVal, comp1744minI, comp1744minJ);
    wire [11:0] comp1745minVal;
    wire [5:0] comp1745minI, comp1745minJ;
    Comparator comp1745(SADValues[3879*12 +: 12], 60, 39, SADValues[3880*12 +: 12], 60, 40, comp1745minVal, comp1745minI, comp1745minJ);
    wire [11:0] comp1746minVal;
    wire [5:0] comp1746minI, comp1746minJ;
    Comparator comp1746(SADValues[3817*12 +: 12], 59, 41, SADValues[3754*12 +: 12], 58, 42, comp1746minVal, comp1746minI, comp1746minJ);
    wire [11:0] comp1747minVal;
    wire [5:0] comp1747minI, comp1747minJ;
    Comparator comp1747(SADValues[3691*12 +: 12], 57, 43, SADValues[3628*12 +: 12], 56, 44, comp1747minVal, comp1747minI, comp1747minJ);
    wire [11:0] comp1748minVal;
    wire [5:0] comp1748minI, comp1748minJ;
    Comparator comp1748(SADValues[3565*12 +: 12], 55, 45, SADValues[3502*12 +: 12], 54, 46, comp1748minVal, comp1748minI, comp1748minJ);
    wire [11:0] comp1749minVal;
    wire [5:0] comp1749minI, comp1749minJ;
    Comparator comp1749(SADValues[3439*12 +: 12], 53, 47, SADValues[3376*12 +: 12], 52, 48, comp1749minVal, comp1749minI, comp1749minJ);
    wire [11:0] comp1750minVal;
    wire [5:0] comp1750minI, comp1750minJ;
    Comparator comp1750(SADValues[3313*12 +: 12], 51, 49, SADValues[3250*12 +: 12], 50, 50, comp1750minVal, comp1750minI, comp1750minJ);
    wire [11:0] comp1751minVal;
    wire [5:0] comp1751minI, comp1751minJ;
    Comparator comp1751(SADValues[3187*12 +: 12], 49, 51, SADValues[3124*12 +: 12], 48, 52, comp1751minVal, comp1751minI, comp1751minJ);
    wire [11:0] comp1752minVal;
    wire [5:0] comp1752minI, comp1752minJ;
    Comparator comp1752(SADValues[3061*12 +: 12], 47, 53, SADValues[2998*12 +: 12], 46, 54, comp1752minVal, comp1752minI, comp1752minJ);
    wire [11:0] comp1753minVal;
    wire [5:0] comp1753minI, comp1753minJ;
    Comparator comp1753(SADValues[2935*12 +: 12], 45, 55, SADValues[2872*12 +: 12], 44, 56, comp1753minVal, comp1753minI, comp1753minJ);
    wire [11:0] comp1754minVal;
    wire [5:0] comp1754minI, comp1754minJ;
    Comparator comp1754(SADValues[2809*12 +: 12], 43, 57, SADValues[2746*12 +: 12], 42, 58, comp1754minVal, comp1754minI, comp1754minJ);
    wire [11:0] comp1755minVal;
    wire [5:0] comp1755minI, comp1755minJ;
    Comparator comp1755(SADValues[2683*12 +: 12], 41, 59, SADValues[2620*12 +: 12], 40, 60, comp1755minVal, comp1755minI, comp1755minJ);
    wire [11:0] comp1756minVal;
    wire [5:0] comp1756minI, comp1756minJ;
    Comparator comp1756(SADValues[2684*12 +: 12], 41, 60, SADValues[2747*12 +: 12], 42, 59, comp1756minVal, comp1756minI, comp1756minJ);
    wire [11:0] comp1757minVal;
    wire [5:0] comp1757minI, comp1757minJ;
    Comparator comp1757(SADValues[2810*12 +: 12], 43, 58, SADValues[2873*12 +: 12], 44, 57, comp1757minVal, comp1757minI, comp1757minJ);
    wire [11:0] comp1758minVal;
    wire [5:0] comp1758minI, comp1758minJ;
    Comparator comp1758(SADValues[2936*12 +: 12], 45, 56, SADValues[2999*12 +: 12], 46, 55, comp1758minVal, comp1758minI, comp1758minJ);
    wire [11:0] comp1759minVal;
    wire [5:0] comp1759minI, comp1759minJ;
    Comparator comp1759(SADValues[3062*12 +: 12], 47, 54, SADValues[3125*12 +: 12], 48, 53, comp1759minVal, comp1759minI, comp1759minJ);
    wire [11:0] comp1760minVal;
    wire [5:0] comp1760minI, comp1760minJ;
    Comparator comp1760(SADValues[3188*12 +: 12], 49, 52, SADValues[3251*12 +: 12], 50, 51, comp1760minVal, comp1760minI, comp1760minJ);
    wire [11:0] comp1761minVal;
    wire [5:0] comp1761minI, comp1761minJ;
    Comparator comp1761(SADValues[3314*12 +: 12], 51, 50, SADValues[3377*12 +: 12], 52, 49, comp1761minVal, comp1761minI, comp1761minJ);
    wire [11:0] comp1762minVal;
    wire [5:0] comp1762minI, comp1762minJ;
    Comparator comp1762(SADValues[3440*12 +: 12], 53, 48, SADValues[3503*12 +: 12], 54, 47, comp1762minVal, comp1762minI, comp1762minJ);
    wire [11:0] comp1763minVal;
    wire [5:0] comp1763minI, comp1763minJ;
    Comparator comp1763(SADValues[3566*12 +: 12], 55, 46, SADValues[3629*12 +: 12], 56, 45, comp1763minVal, comp1763minI, comp1763minJ);
    wire [11:0] comp1764minVal;
    wire [5:0] comp1764minI, comp1764minJ;
    Comparator comp1764(SADValues[3692*12 +: 12], 57, 44, SADValues[3755*12 +: 12], 58, 43, comp1764minVal, comp1764minI, comp1764minJ);
    wire [11:0] comp1765minVal;
    wire [5:0] comp1765minI, comp1765minJ;
    Comparator comp1765(SADValues[3818*12 +: 12], 59, 42, SADValues[3881*12 +: 12], 60, 41, comp1765minVal, comp1765minI, comp1765minJ);
    wire [11:0] comp1766minVal;
    wire [5:0] comp1766minI, comp1766minJ;
    Comparator comp1766(SADValues[3882*12 +: 12], 60, 42, SADValues[3819*12 +: 12], 59, 43, comp1766minVal, comp1766minI, comp1766minJ);
    wire [11:0] comp1767minVal;
    wire [5:0] comp1767minI, comp1767minJ;
    Comparator comp1767(SADValues[3756*12 +: 12], 58, 44, SADValues[3693*12 +: 12], 57, 45, comp1767minVal, comp1767minI, comp1767minJ);
    wire [11:0] comp1768minVal;
    wire [5:0] comp1768minI, comp1768minJ;
    Comparator comp1768(SADValues[3630*12 +: 12], 56, 46, SADValues[3567*12 +: 12], 55, 47, comp1768minVal, comp1768minI, comp1768minJ);
    wire [11:0] comp1769minVal;
    wire [5:0] comp1769minI, comp1769minJ;
    Comparator comp1769(SADValues[3504*12 +: 12], 54, 48, SADValues[3441*12 +: 12], 53, 49, comp1769minVal, comp1769minI, comp1769minJ);
    wire [11:0] comp1770minVal;
    wire [5:0] comp1770minI, comp1770minJ;
    Comparator comp1770(SADValues[3378*12 +: 12], 52, 50, SADValues[3315*12 +: 12], 51, 51, comp1770minVal, comp1770minI, comp1770minJ);
    wire [11:0] comp1771minVal;
    wire [5:0] comp1771minI, comp1771minJ;
    Comparator comp1771(SADValues[3252*12 +: 12], 50, 52, SADValues[3189*12 +: 12], 49, 53, comp1771minVal, comp1771minI, comp1771minJ);
    wire [11:0] comp1772minVal;
    wire [5:0] comp1772minI, comp1772minJ;
    Comparator comp1772(SADValues[3126*12 +: 12], 48, 54, SADValues[3063*12 +: 12], 47, 55, comp1772minVal, comp1772minI, comp1772minJ);
    wire [11:0] comp1773minVal;
    wire [5:0] comp1773minI, comp1773minJ;
    Comparator comp1773(SADValues[3000*12 +: 12], 46, 56, SADValues[2937*12 +: 12], 45, 57, comp1773minVal, comp1773minI, comp1773minJ);
    wire [11:0] comp1774minVal;
    wire [5:0] comp1774minI, comp1774minJ;
    Comparator comp1774(SADValues[2874*12 +: 12], 44, 58, SADValues[2811*12 +: 12], 43, 59, comp1774minVal, comp1774minI, comp1774minJ);
    wire [11:0] comp1775minVal;
    wire [5:0] comp1775minI, comp1775minJ;
    Comparator comp1775(SADValues[2748*12 +: 12], 42, 60, SADValues[2812*12 +: 12], 43, 60, comp1775minVal, comp1775minI, comp1775minJ);
    wire [11:0] comp1776minVal;
    wire [5:0] comp1776minI, comp1776minJ;
    Comparator comp1776(SADValues[2875*12 +: 12], 44, 59, SADValues[2938*12 +: 12], 45, 58, comp1776minVal, comp1776minI, comp1776minJ);
    wire [11:0] comp1777minVal;
    wire [5:0] comp1777minI, comp1777minJ;
    Comparator comp1777(SADValues[3001*12 +: 12], 46, 57, SADValues[3064*12 +: 12], 47, 56, comp1777minVal, comp1777minI, comp1777minJ);
    wire [11:0] comp1778minVal;
    wire [5:0] comp1778minI, comp1778minJ;
    Comparator comp1778(SADValues[3127*12 +: 12], 48, 55, SADValues[3190*12 +: 12], 49, 54, comp1778minVal, comp1778minI, comp1778minJ);
    wire [11:0] comp1779minVal;
    wire [5:0] comp1779minI, comp1779minJ;
    Comparator comp1779(SADValues[3253*12 +: 12], 50, 53, SADValues[3316*12 +: 12], 51, 52, comp1779minVal, comp1779minI, comp1779minJ);
    wire [11:0] comp1780minVal;
    wire [5:0] comp1780minI, comp1780minJ;
    Comparator comp1780(SADValues[3379*12 +: 12], 52, 51, SADValues[3442*12 +: 12], 53, 50, comp1780minVal, comp1780minI, comp1780minJ);
    wire [11:0] comp1781minVal;
    wire [5:0] comp1781minI, comp1781minJ;
    Comparator comp1781(SADValues[3505*12 +: 12], 54, 49, SADValues[3568*12 +: 12], 55, 48, comp1781minVal, comp1781minI, comp1781minJ);
    wire [11:0] comp1782minVal;
    wire [5:0] comp1782minI, comp1782minJ;
    Comparator comp1782(SADValues[3631*12 +: 12], 56, 47, SADValues[3694*12 +: 12], 57, 46, comp1782minVal, comp1782minI, comp1782minJ);
    wire [11:0] comp1783minVal;
    wire [5:0] comp1783minI, comp1783minJ;
    Comparator comp1783(SADValues[3757*12 +: 12], 58, 45, SADValues[3820*12 +: 12], 59, 44, comp1783minVal, comp1783minI, comp1783minJ);
    wire [11:0] comp1784minVal;
    wire [5:0] comp1784minI, comp1784minJ;
    Comparator comp1784(SADValues[3883*12 +: 12], 60, 43, SADValues[3884*12 +: 12], 60, 44, comp1784minVal, comp1784minI, comp1784minJ);
    wire [11:0] comp1785minVal;
    wire [5:0] comp1785minI, comp1785minJ;
    Comparator comp1785(SADValues[3821*12 +: 12], 59, 45, SADValues[3758*12 +: 12], 58, 46, comp1785minVal, comp1785minI, comp1785minJ);
    wire [11:0] comp1786minVal;
    wire [5:0] comp1786minI, comp1786minJ;
    Comparator comp1786(SADValues[3695*12 +: 12], 57, 47, SADValues[3632*12 +: 12], 56, 48, comp1786minVal, comp1786minI, comp1786minJ);
    wire [11:0] comp1787minVal;
    wire [5:0] comp1787minI, comp1787minJ;
    Comparator comp1787(SADValues[3569*12 +: 12], 55, 49, SADValues[3506*12 +: 12], 54, 50, comp1787minVal, comp1787minI, comp1787minJ);
    wire [11:0] comp1788minVal;
    wire [5:0] comp1788minI, comp1788minJ;
    Comparator comp1788(SADValues[3443*12 +: 12], 53, 51, SADValues[3380*12 +: 12], 52, 52, comp1788minVal, comp1788minI, comp1788minJ);
    wire [11:0] comp1789minVal;
    wire [5:0] comp1789minI, comp1789minJ;
    Comparator comp1789(SADValues[3317*12 +: 12], 51, 53, SADValues[3254*12 +: 12], 50, 54, comp1789minVal, comp1789minI, comp1789minJ);
    wire [11:0] comp1790minVal;
    wire [5:0] comp1790minI, comp1790minJ;
    Comparator comp1790(SADValues[3191*12 +: 12], 49, 55, SADValues[3128*12 +: 12], 48, 56, comp1790minVal, comp1790minI, comp1790minJ);
    wire [11:0] comp1791minVal;
    wire [5:0] comp1791minI, comp1791minJ;
    Comparator comp1791(SADValues[3065*12 +: 12], 47, 57, SADValues[3002*12 +: 12], 46, 58, comp1791minVal, comp1791minI, comp1791minJ);
    wire [11:0] comp1792minVal;
    wire [5:0] comp1792minI, comp1792minJ;
    Comparator comp1792(SADValues[2939*12 +: 12], 45, 59, SADValues[2876*12 +: 12], 44, 60, comp1792minVal, comp1792minI, comp1792minJ);
    wire [11:0] comp1793minVal;
    wire [5:0] comp1793minI, comp1793minJ;
    Comparator comp1793(SADValues[2940*12 +: 12], 45, 60, SADValues[3003*12 +: 12], 46, 59, comp1793minVal, comp1793minI, comp1793minJ);
    wire [11:0] comp1794minVal;
    wire [5:0] comp1794minI, comp1794minJ;
    Comparator comp1794(SADValues[3066*12 +: 12], 47, 58, SADValues[3129*12 +: 12], 48, 57, comp1794minVal, comp1794minI, comp1794minJ);
    wire [11:0] comp1795minVal;
    wire [5:0] comp1795minI, comp1795minJ;
    Comparator comp1795(SADValues[3192*12 +: 12], 49, 56, SADValues[3255*12 +: 12], 50, 55, comp1795minVal, comp1795minI, comp1795minJ);
    wire [11:0] comp1796minVal;
    wire [5:0] comp1796minI, comp1796minJ;
    Comparator comp1796(SADValues[3318*12 +: 12], 51, 54, SADValues[3381*12 +: 12], 52, 53, comp1796minVal, comp1796minI, comp1796minJ);
    wire [11:0] comp1797minVal;
    wire [5:0] comp1797minI, comp1797minJ;
    Comparator comp1797(SADValues[3444*12 +: 12], 53, 52, SADValues[3507*12 +: 12], 54, 51, comp1797minVal, comp1797minI, comp1797minJ);
    wire [11:0] comp1798minVal;
    wire [5:0] comp1798minI, comp1798minJ;
    Comparator comp1798(SADValues[3570*12 +: 12], 55, 50, SADValues[3633*12 +: 12], 56, 49, comp1798minVal, comp1798minI, comp1798minJ);
    wire [11:0] comp1799minVal;
    wire [5:0] comp1799minI, comp1799minJ;
    Comparator comp1799(SADValues[3696*12 +: 12], 57, 48, SADValues[3759*12 +: 12], 58, 47, comp1799minVal, comp1799minI, comp1799minJ);
    wire [11:0] comp1800minVal;
    wire [5:0] comp1800minI, comp1800minJ;
    Comparator comp1800(SADValues[3822*12 +: 12], 59, 46, SADValues[3885*12 +: 12], 60, 45, comp1800minVal, comp1800minI, comp1800minJ);
    wire [11:0] comp1801minVal;
    wire [5:0] comp1801minI, comp1801minJ;
    Comparator comp1801(SADValues[3886*12 +: 12], 60, 46, SADValues[3823*12 +: 12], 59, 47, comp1801minVal, comp1801minI, comp1801minJ);
    wire [11:0] comp1802minVal;
    wire [5:0] comp1802minI, comp1802minJ;
    Comparator comp1802(SADValues[3760*12 +: 12], 58, 48, SADValues[3697*12 +: 12], 57, 49, comp1802minVal, comp1802minI, comp1802minJ);
    wire [11:0] comp1803minVal;
    wire [5:0] comp1803minI, comp1803minJ;
    Comparator comp1803(SADValues[3634*12 +: 12], 56, 50, SADValues[3571*12 +: 12], 55, 51, comp1803minVal, comp1803minI, comp1803minJ);
    wire [11:0] comp1804minVal;
    wire [5:0] comp1804minI, comp1804minJ;
    Comparator comp1804(SADValues[3508*12 +: 12], 54, 52, SADValues[3445*12 +: 12], 53, 53, comp1804minVal, comp1804minI, comp1804minJ);
    wire [11:0] comp1805minVal;
    wire [5:0] comp1805minI, comp1805minJ;
    Comparator comp1805(SADValues[3382*12 +: 12], 52, 54, SADValues[3319*12 +: 12], 51, 55, comp1805minVal, comp1805minI, comp1805minJ);
    wire [11:0] comp1806minVal;
    wire [5:0] comp1806minI, comp1806minJ;
    Comparator comp1806(SADValues[3256*12 +: 12], 50, 56, SADValues[3193*12 +: 12], 49, 57, comp1806minVal, comp1806minI, comp1806minJ);
    wire [11:0] comp1807minVal;
    wire [5:0] comp1807minI, comp1807minJ;
    Comparator comp1807(SADValues[3130*12 +: 12], 48, 58, SADValues[3067*12 +: 12], 47, 59, comp1807minVal, comp1807minI, comp1807minJ);
    wire [11:0] comp1808minVal;
    wire [5:0] comp1808minI, comp1808minJ;
    Comparator comp1808(SADValues[3004*12 +: 12], 46, 60, SADValues[3068*12 +: 12], 47, 60, comp1808minVal, comp1808minI, comp1808minJ);
    wire [11:0] comp1809minVal;
    wire [5:0] comp1809minI, comp1809minJ;
    Comparator comp1809(SADValues[3131*12 +: 12], 48, 59, SADValues[3194*12 +: 12], 49, 58, comp1809minVal, comp1809minI, comp1809minJ);
    wire [11:0] comp1810minVal;
    wire [5:0] comp1810minI, comp1810minJ;
    Comparator comp1810(SADValues[3257*12 +: 12], 50, 57, SADValues[3320*12 +: 12], 51, 56, comp1810minVal, comp1810minI, comp1810minJ);
    wire [11:0] comp1811minVal;
    wire [5:0] comp1811minI, comp1811minJ;
    Comparator comp1811(SADValues[3383*12 +: 12], 52, 55, SADValues[3446*12 +: 12], 53, 54, comp1811minVal, comp1811minI, comp1811minJ);
    wire [11:0] comp1812minVal;
    wire [5:0] comp1812minI, comp1812minJ;
    Comparator comp1812(SADValues[3509*12 +: 12], 54, 53, SADValues[3572*12 +: 12], 55, 52, comp1812minVal, comp1812minI, comp1812minJ);
    wire [11:0] comp1813minVal;
    wire [5:0] comp1813minI, comp1813minJ;
    Comparator comp1813(SADValues[3635*12 +: 12], 56, 51, SADValues[3698*12 +: 12], 57, 50, comp1813minVal, comp1813minI, comp1813minJ);
    wire [11:0] comp1814minVal;
    wire [5:0] comp1814minI, comp1814minJ;
    Comparator comp1814(SADValues[3761*12 +: 12], 58, 49, SADValues[3824*12 +: 12], 59, 48, comp1814minVal, comp1814minI, comp1814minJ);
    wire [11:0] comp1815minVal;
    wire [5:0] comp1815minI, comp1815minJ;
    Comparator comp1815(SADValues[3887*12 +: 12], 60, 47, SADValues[3888*12 +: 12], 60, 48, comp1815minVal, comp1815minI, comp1815minJ);
    wire [11:0] comp1816minVal;
    wire [5:0] comp1816minI, comp1816minJ;
    Comparator comp1816(SADValues[3825*12 +: 12], 59, 49, SADValues[3762*12 +: 12], 58, 50, comp1816minVal, comp1816minI, comp1816minJ);
    wire [11:0] comp1817minVal;
    wire [5:0] comp1817minI, comp1817minJ;
    Comparator comp1817(SADValues[3699*12 +: 12], 57, 51, SADValues[3636*12 +: 12], 56, 52, comp1817minVal, comp1817minI, comp1817minJ);
    wire [11:0] comp1818minVal;
    wire [5:0] comp1818minI, comp1818minJ;
    Comparator comp1818(SADValues[3573*12 +: 12], 55, 53, SADValues[3510*12 +: 12], 54, 54, comp1818minVal, comp1818minI, comp1818minJ);
    wire [11:0] comp1819minVal;
    wire [5:0] comp1819minI, comp1819minJ;
    Comparator comp1819(SADValues[3447*12 +: 12], 53, 55, SADValues[3384*12 +: 12], 52, 56, comp1819minVal, comp1819minI, comp1819minJ);
    wire [11:0] comp1820minVal;
    wire [5:0] comp1820minI, comp1820minJ;
    Comparator comp1820(SADValues[3321*12 +: 12], 51, 57, SADValues[3258*12 +: 12], 50, 58, comp1820minVal, comp1820minI, comp1820minJ);
    wire [11:0] comp1821minVal;
    wire [5:0] comp1821minI, comp1821minJ;
    Comparator comp1821(SADValues[3195*12 +: 12], 49, 59, SADValues[3132*12 +: 12], 48, 60, comp1821minVal, comp1821minI, comp1821minJ);
    wire [11:0] comp1822minVal;
    wire [5:0] comp1822minI, comp1822minJ;
    Comparator comp1822(SADValues[3196*12 +: 12], 49, 60, SADValues[3259*12 +: 12], 50, 59, comp1822minVal, comp1822minI, comp1822minJ);
    wire [11:0] comp1823minVal;
    wire [5:0] comp1823minI, comp1823minJ;
    Comparator comp1823(SADValues[3322*12 +: 12], 51, 58, SADValues[3385*12 +: 12], 52, 57, comp1823minVal, comp1823minI, comp1823minJ);
    wire [11:0] comp1824minVal;
    wire [5:0] comp1824minI, comp1824minJ;
    Comparator comp1824(SADValues[3448*12 +: 12], 53, 56, SADValues[3511*12 +: 12], 54, 55, comp1824minVal, comp1824minI, comp1824minJ);
    wire [11:0] comp1825minVal;
    wire [5:0] comp1825minI, comp1825minJ;
    Comparator comp1825(SADValues[3574*12 +: 12], 55, 54, SADValues[3637*12 +: 12], 56, 53, comp1825minVal, comp1825minI, comp1825minJ);
    wire [11:0] comp1826minVal;
    wire [5:0] comp1826minI, comp1826minJ;
    Comparator comp1826(SADValues[3700*12 +: 12], 57, 52, SADValues[3763*12 +: 12], 58, 51, comp1826minVal, comp1826minI, comp1826minJ);
    wire [11:0] comp1827minVal;
    wire [5:0] comp1827minI, comp1827minJ;
    Comparator comp1827(SADValues[3826*12 +: 12], 59, 50, SADValues[3889*12 +: 12], 60, 49, comp1827minVal, comp1827minI, comp1827minJ);
    wire [11:0] comp1828minVal;
    wire [5:0] comp1828minI, comp1828minJ;
    Comparator comp1828(SADValues[3890*12 +: 12], 60, 50, SADValues[3827*12 +: 12], 59, 51, comp1828minVal, comp1828minI, comp1828minJ);
    wire [11:0] comp1829minVal;
    wire [5:0] comp1829minI, comp1829minJ;
    Comparator comp1829(SADValues[3764*12 +: 12], 58, 52, SADValues[3701*12 +: 12], 57, 53, comp1829minVal, comp1829minI, comp1829minJ);
    wire [11:0] comp1830minVal;
    wire [5:0] comp1830minI, comp1830minJ;
    Comparator comp1830(SADValues[3638*12 +: 12], 56, 54, SADValues[3575*12 +: 12], 55, 55, comp1830minVal, comp1830minI, comp1830minJ);
    wire [11:0] comp1831minVal;
    wire [5:0] comp1831minI, comp1831minJ;
    Comparator comp1831(SADValues[3512*12 +: 12], 54, 56, SADValues[3449*12 +: 12], 53, 57, comp1831minVal, comp1831minI, comp1831minJ);
    wire [11:0] comp1832minVal;
    wire [5:0] comp1832minI, comp1832minJ;
    Comparator comp1832(SADValues[3386*12 +: 12], 52, 58, SADValues[3323*12 +: 12], 51, 59, comp1832minVal, comp1832minI, comp1832minJ);
    wire [11:0] comp1833minVal;
    wire [5:0] comp1833minI, comp1833minJ;
    Comparator comp1833(SADValues[3260*12 +: 12], 50, 60, SADValues[3324*12 +: 12], 51, 60, comp1833minVal, comp1833minI, comp1833minJ);
    wire [11:0] comp1834minVal;
    wire [5:0] comp1834minI, comp1834minJ;
    Comparator comp1834(SADValues[3387*12 +: 12], 52, 59, SADValues[3450*12 +: 12], 53, 58, comp1834minVal, comp1834minI, comp1834minJ);
    wire [11:0] comp1835minVal;
    wire [5:0] comp1835minI, comp1835minJ;
    Comparator comp1835(SADValues[3513*12 +: 12], 54, 57, SADValues[3576*12 +: 12], 55, 56, comp1835minVal, comp1835minI, comp1835minJ);
    wire [11:0] comp1836minVal;
    wire [5:0] comp1836minI, comp1836minJ;
    Comparator comp1836(SADValues[3639*12 +: 12], 56, 55, SADValues[3702*12 +: 12], 57, 54, comp1836minVal, comp1836minI, comp1836minJ);
    wire [11:0] comp1837minVal;
    wire [5:0] comp1837minI, comp1837minJ;
    Comparator comp1837(SADValues[3765*12 +: 12], 58, 53, SADValues[3828*12 +: 12], 59, 52, comp1837minVal, comp1837minI, comp1837minJ);
    wire [11:0] comp1838minVal;
    wire [5:0] comp1838minI, comp1838minJ;
    Comparator comp1838(SADValues[3891*12 +: 12], 60, 51, SADValues[3892*12 +: 12], 60, 52, comp1838minVal, comp1838minI, comp1838minJ);
    wire [11:0] comp1839minVal;
    wire [5:0] comp1839minI, comp1839minJ;
    Comparator comp1839(SADValues[3829*12 +: 12], 59, 53, SADValues[3766*12 +: 12], 58, 54, comp1839minVal, comp1839minI, comp1839minJ);
    wire [11:0] comp1840minVal;
    wire [5:0] comp1840minI, comp1840minJ;
    Comparator comp1840(SADValues[3703*12 +: 12], 57, 55, SADValues[3640*12 +: 12], 56, 56, comp1840minVal, comp1840minI, comp1840minJ);
    wire [11:0] comp1841minVal;
    wire [5:0] comp1841minI, comp1841minJ;
    Comparator comp1841(SADValues[3577*12 +: 12], 55, 57, SADValues[3514*12 +: 12], 54, 58, comp1841minVal, comp1841minI, comp1841minJ);
    wire [11:0] comp1842minVal;
    wire [5:0] comp1842minI, comp1842minJ;
    Comparator comp1842(SADValues[3451*12 +: 12], 53, 59, SADValues[3388*12 +: 12], 52, 60, comp1842minVal, comp1842minI, comp1842minJ);
    wire [11:0] comp1843minVal;
    wire [5:0] comp1843minI, comp1843minJ;
    Comparator comp1843(SADValues[3452*12 +: 12], 53, 60, SADValues[3515*12 +: 12], 54, 59, comp1843minVal, comp1843minI, comp1843minJ);
    wire [11:0] comp1844minVal;
    wire [5:0] comp1844minI, comp1844minJ;
    Comparator comp1844(SADValues[3578*12 +: 12], 55, 58, SADValues[3641*12 +: 12], 56, 57, comp1844minVal, comp1844minI, comp1844minJ);
    wire [11:0] comp1845minVal;
    wire [5:0] comp1845minI, comp1845minJ;
    Comparator comp1845(SADValues[3704*12 +: 12], 57, 56, SADValues[3767*12 +: 12], 58, 55, comp1845minVal, comp1845minI, comp1845minJ);
    wire [11:0] comp1846minVal;
    wire [5:0] comp1846minI, comp1846minJ;
    Comparator comp1846(SADValues[3830*12 +: 12], 59, 54, SADValues[3893*12 +: 12], 60, 53, comp1846minVal, comp1846minI, comp1846minJ);
    wire [11:0] comp1847minVal;
    wire [5:0] comp1847minI, comp1847minJ;
    Comparator comp1847(SADValues[3894*12 +: 12], 60, 54, SADValues[3831*12 +: 12], 59, 55, comp1847minVal, comp1847minI, comp1847minJ);
    wire [11:0] comp1848minVal;
    wire [5:0] comp1848minI, comp1848minJ;
    Comparator comp1848(SADValues[3768*12 +: 12], 58, 56, SADValues[3705*12 +: 12], 57, 57, comp1848minVal, comp1848minI, comp1848minJ);
    wire [11:0] comp1849minVal;
    wire [5:0] comp1849minI, comp1849minJ;
    Comparator comp1849(SADValues[3642*12 +: 12], 56, 58, SADValues[3579*12 +: 12], 55, 59, comp1849minVal, comp1849minI, comp1849minJ);
    wire [11:0] comp1850minVal;
    wire [5:0] comp1850minI, comp1850minJ;
    Comparator comp1850(SADValues[3516*12 +: 12], 54, 60, SADValues[3580*12 +: 12], 55, 60, comp1850minVal, comp1850minI, comp1850minJ);
    wire [11:0] comp1851minVal;
    wire [5:0] comp1851minI, comp1851minJ;
    Comparator comp1851(SADValues[3643*12 +: 12], 56, 59, SADValues[3706*12 +: 12], 57, 58, comp1851minVal, comp1851minI, comp1851minJ);
    wire [11:0] comp1852minVal;
    wire [5:0] comp1852minI, comp1852minJ;
    Comparator comp1852(SADValues[3769*12 +: 12], 58, 57, SADValues[3832*12 +: 12], 59, 56, comp1852minVal, comp1852minI, comp1852minJ);
    wire [11:0] comp1853minVal;
    wire [5:0] comp1853minI, comp1853minJ;
    Comparator comp1853(SADValues[3895*12 +: 12], 60, 55, SADValues[3896*12 +: 12], 60, 56, comp1853minVal, comp1853minI, comp1853minJ);
    wire [11:0] comp1854minVal;
    wire [5:0] comp1854minI, comp1854minJ;
    Comparator comp1854(SADValues[3833*12 +: 12], 59, 57, SADValues[3770*12 +: 12], 58, 58, comp1854minVal, comp1854minI, comp1854minJ);
    wire [11:0] comp1855minVal;
    wire [5:0] comp1855minI, comp1855minJ;
    Comparator comp1855(SADValues[3707*12 +: 12], 57, 59, SADValues[3644*12 +: 12], 56, 60, comp1855minVal, comp1855minI, comp1855minJ);
    wire [11:0] comp1856minVal;
    wire [5:0] comp1856minI, comp1856minJ;
    Comparator comp1856(SADValues[3708*12 +: 12], 57, 60, SADValues[3771*12 +: 12], 58, 59, comp1856minVal, comp1856minI, comp1856minJ);
    wire [11:0] comp1857minVal;
    wire [5:0] comp1857minI, comp1857minJ;
    Comparator comp1857(SADValues[3834*12 +: 12], 59, 58, SADValues[3897*12 +: 12], 60, 57, comp1857minVal, comp1857minI, comp1857minJ);
    wire [11:0] comp1858minVal;
    wire [5:0] comp1858minI, comp1858minJ;
    Comparator comp1858(SADValues[3898*12 +: 12], 60, 58, SADValues[3835*12 +: 12], 59, 59, comp1858minVal, comp1858minI, comp1858minJ);
    wire [11:0] comp1859minVal;
    wire [5:0] comp1859minI, comp1859minJ;
    Comparator comp1859(SADValues[3772*12 +: 12], 58, 60, SADValues[3836*12 +: 12], 59, 60, comp1859minVal, comp1859minI, comp1859minJ);
    wire [11:0] comp1860minVal;
    wire [5:0] comp1860minI, comp1860minJ;
    Comparator comp1860(SADValues[3899*12 +: 12], 60, 59, SADValues[3900*12 +: 12], 60, 60, comp1860minVal, comp1860minI, comp1860minJ);
    wire [11:0] comp1861minVal;
    wire [5:0] comp1861minI, comp1861minJ;
    assign comp1861minVal = 4095;
    assign comp1861minI = 0;
    assign comp1861minJ = 0;
    wire [11:0] comp1862minVal;
    wire [5:0] comp1862minI, comp1862minJ;
    Comparator comp1862(comp0minVal, comp0minI, comp0minJ, comp1minVal, comp1minI, comp1minJ, comp1862minVal, comp1862minI, comp1862minJ);
    wire [11:0] comp1863minVal;
    wire [5:0] comp1863minI, comp1863minJ;
    Comparator comp1863(comp2minVal, comp2minI, comp2minJ, comp3minVal, comp3minI, comp3minJ, comp1863minVal, comp1863minI, comp1863minJ);
    wire [11:0] comp1864minVal;
    wire [5:0] comp1864minI, comp1864minJ;
    Comparator comp1864(comp4minVal, comp4minI, comp4minJ, comp5minVal, comp5minI, comp5minJ, comp1864minVal, comp1864minI, comp1864minJ);
    wire [11:0] comp1865minVal;
    wire [5:0] comp1865minI, comp1865minJ;
    Comparator comp1865(comp6minVal, comp6minI, comp6minJ, comp7minVal, comp7minI, comp7minJ, comp1865minVal, comp1865minI, comp1865minJ);
    wire [11:0] comp1866minVal;
    wire [5:0] comp1866minI, comp1866minJ;
    Comparator comp1866(comp8minVal, comp8minI, comp8minJ, comp9minVal, comp9minI, comp9minJ, comp1866minVal, comp1866minI, comp1866minJ);
    wire [11:0] comp1867minVal;
    wire [5:0] comp1867minI, comp1867minJ;
    Comparator comp1867(comp10minVal, comp10minI, comp10minJ, comp11minVal, comp11minI, comp11minJ, comp1867minVal, comp1867minI, comp1867minJ);
    wire [11:0] comp1868minVal;
    wire [5:0] comp1868minI, comp1868minJ;
    Comparator comp1868(comp12minVal, comp12minI, comp12minJ, comp13minVal, comp13minI, comp13minJ, comp1868minVal, comp1868minI, comp1868minJ);
    wire [11:0] comp1869minVal;
    wire [5:0] comp1869minI, comp1869minJ;
    Comparator comp1869(comp14minVal, comp14minI, comp14minJ, comp15minVal, comp15minI, comp15minJ, comp1869minVal, comp1869minI, comp1869minJ);
    wire [11:0] comp1870minVal;
    wire [5:0] comp1870minI, comp1870minJ;
    Comparator comp1870(comp16minVal, comp16minI, comp16minJ, comp17minVal, comp17minI, comp17minJ, comp1870minVal, comp1870minI, comp1870minJ);
    wire [11:0] comp1871minVal;
    wire [5:0] comp1871minI, comp1871minJ;
    Comparator comp1871(comp18minVal, comp18minI, comp18minJ, comp19minVal, comp19minI, comp19minJ, comp1871minVal, comp1871minI, comp1871minJ);
    wire [11:0] comp1872minVal;
    wire [5:0] comp1872minI, comp1872minJ;
    Comparator comp1872(comp20minVal, comp20minI, comp20minJ, comp21minVal, comp21minI, comp21minJ, comp1872minVal, comp1872minI, comp1872minJ);
    wire [11:0] comp1873minVal;
    wire [5:0] comp1873minI, comp1873minJ;
    Comparator comp1873(comp22minVal, comp22minI, comp22minJ, comp23minVal, comp23minI, comp23minJ, comp1873minVal, comp1873minI, comp1873minJ);
    wire [11:0] comp1874minVal;
    wire [5:0] comp1874minI, comp1874minJ;
    Comparator comp1874(comp24minVal, comp24minI, comp24minJ, comp25minVal, comp25minI, comp25minJ, comp1874minVal, comp1874minI, comp1874minJ);
    wire [11:0] comp1875minVal;
    wire [5:0] comp1875minI, comp1875minJ;
    Comparator comp1875(comp26minVal, comp26minI, comp26minJ, comp27minVal, comp27minI, comp27minJ, comp1875minVal, comp1875minI, comp1875minJ);
    wire [11:0] comp1876minVal;
    wire [5:0] comp1876minI, comp1876minJ;
    Comparator comp1876(comp28minVal, comp28minI, comp28minJ, comp29minVal, comp29minI, comp29minJ, comp1876minVal, comp1876minI, comp1876minJ);
    wire [11:0] comp1877minVal;
    wire [5:0] comp1877minI, comp1877minJ;
    Comparator comp1877(comp30minVal, comp30minI, comp30minJ, comp31minVal, comp31minI, comp31minJ, comp1877minVal, comp1877minI, comp1877minJ);
    wire [11:0] comp1878minVal;
    wire [5:0] comp1878minI, comp1878minJ;
    Comparator comp1878(comp32minVal, comp32minI, comp32minJ, comp33minVal, comp33minI, comp33minJ, comp1878minVal, comp1878minI, comp1878minJ);
    wire [11:0] comp1879minVal;
    wire [5:0] comp1879minI, comp1879minJ;
    Comparator comp1879(comp34minVal, comp34minI, comp34minJ, comp35minVal, comp35minI, comp35minJ, comp1879minVal, comp1879minI, comp1879minJ);
    wire [11:0] comp1880minVal;
    wire [5:0] comp1880minI, comp1880minJ;
    Comparator comp1880(comp36minVal, comp36minI, comp36minJ, comp37minVal, comp37minI, comp37minJ, comp1880minVal, comp1880minI, comp1880minJ);
    wire [11:0] comp1881minVal;
    wire [5:0] comp1881minI, comp1881minJ;
    Comparator comp1881(comp38minVal, comp38minI, comp38minJ, comp39minVal, comp39minI, comp39minJ, comp1881minVal, comp1881minI, comp1881minJ);
    wire [11:0] comp1882minVal;
    wire [5:0] comp1882minI, comp1882minJ;
    Comparator comp1882(comp40minVal, comp40minI, comp40minJ, comp41minVal, comp41minI, comp41minJ, comp1882minVal, comp1882minI, comp1882minJ);
    wire [11:0] comp1883minVal;
    wire [5:0] comp1883minI, comp1883minJ;
    Comparator comp1883(comp42minVal, comp42minI, comp42minJ, comp43minVal, comp43minI, comp43minJ, comp1883minVal, comp1883minI, comp1883minJ);
    wire [11:0] comp1884minVal;
    wire [5:0] comp1884minI, comp1884minJ;
    Comparator comp1884(comp44minVal, comp44minI, comp44minJ, comp45minVal, comp45minI, comp45minJ, comp1884minVal, comp1884minI, comp1884minJ);
    wire [11:0] comp1885minVal;
    wire [5:0] comp1885minI, comp1885minJ;
    Comparator comp1885(comp46minVal, comp46minI, comp46minJ, comp47minVal, comp47minI, comp47minJ, comp1885minVal, comp1885minI, comp1885minJ);
    wire [11:0] comp1886minVal;
    wire [5:0] comp1886minI, comp1886minJ;
    Comparator comp1886(comp48minVal, comp48minI, comp48minJ, comp49minVal, comp49minI, comp49minJ, comp1886minVal, comp1886minI, comp1886minJ);
    wire [11:0] comp1887minVal;
    wire [5:0] comp1887minI, comp1887minJ;
    Comparator comp1887(comp50minVal, comp50minI, comp50minJ, comp51minVal, comp51minI, comp51minJ, comp1887minVal, comp1887minI, comp1887minJ);
    wire [11:0] comp1888minVal;
    wire [5:0] comp1888minI, comp1888minJ;
    Comparator comp1888(comp52minVal, comp52minI, comp52minJ, comp53minVal, comp53minI, comp53minJ, comp1888minVal, comp1888minI, comp1888minJ);
    wire [11:0] comp1889minVal;
    wire [5:0] comp1889minI, comp1889minJ;
    Comparator comp1889(comp54minVal, comp54minI, comp54minJ, comp55minVal, comp55minI, comp55minJ, comp1889minVal, comp1889minI, comp1889minJ);
    wire [11:0] comp1890minVal;
    wire [5:0] comp1890minI, comp1890minJ;
    Comparator comp1890(comp56minVal, comp56minI, comp56minJ, comp57minVal, comp57minI, comp57minJ, comp1890minVal, comp1890minI, comp1890minJ);
    wire [11:0] comp1891minVal;
    wire [5:0] comp1891minI, comp1891minJ;
    Comparator comp1891(comp58minVal, comp58minI, comp58minJ, comp59minVal, comp59minI, comp59minJ, comp1891minVal, comp1891minI, comp1891minJ);
    wire [11:0] comp1892minVal;
    wire [5:0] comp1892minI, comp1892minJ;
    Comparator comp1892(comp60minVal, comp60minI, comp60minJ, comp61minVal, comp61minI, comp61minJ, comp1892minVal, comp1892minI, comp1892minJ);
    wire [11:0] comp1893minVal;
    wire [5:0] comp1893minI, comp1893minJ;
    Comparator comp1893(comp62minVal, comp62minI, comp62minJ, comp63minVal, comp63minI, comp63minJ, comp1893minVal, comp1893minI, comp1893minJ);
    wire [11:0] comp1894minVal;
    wire [5:0] comp1894minI, comp1894minJ;
    Comparator comp1894(comp64minVal, comp64minI, comp64minJ, comp65minVal, comp65minI, comp65minJ, comp1894minVal, comp1894minI, comp1894minJ);
    wire [11:0] comp1895minVal;
    wire [5:0] comp1895minI, comp1895minJ;
    Comparator comp1895(comp66minVal, comp66minI, comp66minJ, comp67minVal, comp67minI, comp67minJ, comp1895minVal, comp1895minI, comp1895minJ);
    wire [11:0] comp1896minVal;
    wire [5:0] comp1896minI, comp1896minJ;
    Comparator comp1896(comp68minVal, comp68minI, comp68minJ, comp69minVal, comp69minI, comp69minJ, comp1896minVal, comp1896minI, comp1896minJ);
    wire [11:0] comp1897minVal;
    wire [5:0] comp1897minI, comp1897minJ;
    Comparator comp1897(comp70minVal, comp70minI, comp70minJ, comp71minVal, comp71minI, comp71minJ, comp1897minVal, comp1897minI, comp1897minJ);
    wire [11:0] comp1898minVal;
    wire [5:0] comp1898minI, comp1898minJ;
    Comparator comp1898(comp72minVal, comp72minI, comp72minJ, comp73minVal, comp73minI, comp73minJ, comp1898minVal, comp1898minI, comp1898minJ);
    wire [11:0] comp1899minVal;
    wire [5:0] comp1899minI, comp1899minJ;
    Comparator comp1899(comp74minVal, comp74minI, comp74minJ, comp75minVal, comp75minI, comp75minJ, comp1899minVal, comp1899minI, comp1899minJ);
    wire [11:0] comp1900minVal;
    wire [5:0] comp1900minI, comp1900minJ;
    Comparator comp1900(comp76minVal, comp76minI, comp76minJ, comp77minVal, comp77minI, comp77minJ, comp1900minVal, comp1900minI, comp1900minJ);
    wire [11:0] comp1901minVal;
    wire [5:0] comp1901minI, comp1901minJ;
    Comparator comp1901(comp78minVal, comp78minI, comp78minJ, comp79minVal, comp79minI, comp79minJ, comp1901minVal, comp1901minI, comp1901minJ);
    wire [11:0] comp1902minVal;
    wire [5:0] comp1902minI, comp1902minJ;
    Comparator comp1902(comp80minVal, comp80minI, comp80minJ, comp81minVal, comp81minI, comp81minJ, comp1902minVal, comp1902minI, comp1902minJ);
    wire [11:0] comp1903minVal;
    wire [5:0] comp1903minI, comp1903minJ;
    Comparator comp1903(comp82minVal, comp82minI, comp82minJ, comp83minVal, comp83minI, comp83minJ, comp1903minVal, comp1903minI, comp1903minJ);
    wire [11:0] comp1904minVal;
    wire [5:0] comp1904minI, comp1904minJ;
    Comparator comp1904(comp84minVal, comp84minI, comp84minJ, comp85minVal, comp85minI, comp85minJ, comp1904minVal, comp1904minI, comp1904minJ);
    wire [11:0] comp1905minVal;
    wire [5:0] comp1905minI, comp1905minJ;
    Comparator comp1905(comp86minVal, comp86minI, comp86minJ, comp87minVal, comp87minI, comp87minJ, comp1905minVal, comp1905minI, comp1905minJ);
    wire [11:0] comp1906minVal;
    wire [5:0] comp1906minI, comp1906minJ;
    Comparator comp1906(comp88minVal, comp88minI, comp88minJ, comp89minVal, comp89minI, comp89minJ, comp1906minVal, comp1906minI, comp1906minJ);
    wire [11:0] comp1907minVal;
    wire [5:0] comp1907minI, comp1907minJ;
    Comparator comp1907(comp90minVal, comp90minI, comp90minJ, comp91minVal, comp91minI, comp91minJ, comp1907minVal, comp1907minI, comp1907minJ);
    wire [11:0] comp1908minVal;
    wire [5:0] comp1908minI, comp1908minJ;
    Comparator comp1908(comp92minVal, comp92minI, comp92minJ, comp93minVal, comp93minI, comp93minJ, comp1908minVal, comp1908minI, comp1908minJ);
    wire [11:0] comp1909minVal;
    wire [5:0] comp1909minI, comp1909minJ;
    Comparator comp1909(comp94minVal, comp94minI, comp94minJ, comp95minVal, comp95minI, comp95minJ, comp1909minVal, comp1909minI, comp1909minJ);
    wire [11:0] comp1910minVal;
    wire [5:0] comp1910minI, comp1910minJ;
    Comparator comp1910(comp96minVal, comp96minI, comp96minJ, comp97minVal, comp97minI, comp97minJ, comp1910minVal, comp1910minI, comp1910minJ);
    wire [11:0] comp1911minVal;
    wire [5:0] comp1911minI, comp1911minJ;
    Comparator comp1911(comp98minVal, comp98minI, comp98minJ, comp99minVal, comp99minI, comp99minJ, comp1911minVal, comp1911minI, comp1911minJ);
    wire [11:0] comp1912minVal;
    wire [5:0] comp1912minI, comp1912minJ;
    Comparator comp1912(comp100minVal, comp100minI, comp100minJ, comp101minVal, comp101minI, comp101minJ, comp1912minVal, comp1912minI, comp1912minJ);
    wire [11:0] comp1913minVal;
    wire [5:0] comp1913minI, comp1913minJ;
    Comparator comp1913(comp102minVal, comp102minI, comp102minJ, comp103minVal, comp103minI, comp103minJ, comp1913minVal, comp1913minI, comp1913minJ);
    wire [11:0] comp1914minVal;
    wire [5:0] comp1914minI, comp1914minJ;
    Comparator comp1914(comp104minVal, comp104minI, comp104minJ, comp105minVal, comp105minI, comp105minJ, comp1914minVal, comp1914minI, comp1914minJ);
    wire [11:0] comp1915minVal;
    wire [5:0] comp1915minI, comp1915minJ;
    Comparator comp1915(comp106minVal, comp106minI, comp106minJ, comp107minVal, comp107minI, comp107minJ, comp1915minVal, comp1915minI, comp1915minJ);
    wire [11:0] comp1916minVal;
    wire [5:0] comp1916minI, comp1916minJ;
    Comparator comp1916(comp108minVal, comp108minI, comp108minJ, comp109minVal, comp109minI, comp109minJ, comp1916minVal, comp1916minI, comp1916minJ);
    wire [11:0] comp1917minVal;
    wire [5:0] comp1917minI, comp1917minJ;
    Comparator comp1917(comp110minVal, comp110minI, comp110minJ, comp111minVal, comp111minI, comp111minJ, comp1917minVal, comp1917minI, comp1917minJ);
    wire [11:0] comp1918minVal;
    wire [5:0] comp1918minI, comp1918minJ;
    Comparator comp1918(comp112minVal, comp112minI, comp112minJ, comp113minVal, comp113minI, comp113minJ, comp1918minVal, comp1918minI, comp1918minJ);
    wire [11:0] comp1919minVal;
    wire [5:0] comp1919minI, comp1919minJ;
    Comparator comp1919(comp114minVal, comp114minI, comp114minJ, comp115minVal, comp115minI, comp115minJ, comp1919minVal, comp1919minI, comp1919minJ);
    wire [11:0] comp1920minVal;
    wire [5:0] comp1920minI, comp1920minJ;
    Comparator comp1920(comp116minVal, comp116minI, comp116minJ, comp117minVal, comp117minI, comp117minJ, comp1920minVal, comp1920minI, comp1920minJ);
    wire [11:0] comp1921minVal;
    wire [5:0] comp1921minI, comp1921minJ;
    Comparator comp1921(comp118minVal, comp118minI, comp118minJ, comp119minVal, comp119minI, comp119minJ, comp1921minVal, comp1921minI, comp1921minJ);
    wire [11:0] comp1922minVal;
    wire [5:0] comp1922minI, comp1922minJ;
    Comparator comp1922(comp120minVal, comp120minI, comp120minJ, comp121minVal, comp121minI, comp121minJ, comp1922minVal, comp1922minI, comp1922minJ);
    wire [11:0] comp1923minVal;
    wire [5:0] comp1923minI, comp1923minJ;
    Comparator comp1923(comp122minVal, comp122minI, comp122minJ, comp123minVal, comp123minI, comp123minJ, comp1923minVal, comp1923minI, comp1923minJ);
    wire [11:0] comp1924minVal;
    wire [5:0] comp1924minI, comp1924minJ;
    Comparator comp1924(comp124minVal, comp124minI, comp124minJ, comp125minVal, comp125minI, comp125minJ, comp1924minVal, comp1924minI, comp1924minJ);
    wire [11:0] comp1925minVal;
    wire [5:0] comp1925minI, comp1925minJ;
    Comparator comp1925(comp126minVal, comp126minI, comp126minJ, comp127minVal, comp127minI, comp127minJ, comp1925minVal, comp1925minI, comp1925minJ);
    wire [11:0] comp1926minVal;
    wire [5:0] comp1926minI, comp1926minJ;
    Comparator comp1926(comp128minVal, comp128minI, comp128minJ, comp129minVal, comp129minI, comp129minJ, comp1926minVal, comp1926minI, comp1926minJ);
    wire [11:0] comp1927minVal;
    wire [5:0] comp1927minI, comp1927minJ;
    Comparator comp1927(comp130minVal, comp130minI, comp130minJ, comp131minVal, comp131minI, comp131minJ, comp1927minVal, comp1927minI, comp1927minJ);
    wire [11:0] comp1928minVal;
    wire [5:0] comp1928minI, comp1928minJ;
    Comparator comp1928(comp132minVal, comp132minI, comp132minJ, comp133minVal, comp133minI, comp133minJ, comp1928minVal, comp1928minI, comp1928minJ);
    wire [11:0] comp1929minVal;
    wire [5:0] comp1929minI, comp1929minJ;
    Comparator comp1929(comp134minVal, comp134minI, comp134minJ, comp135minVal, comp135minI, comp135minJ, comp1929minVal, comp1929minI, comp1929minJ);
    wire [11:0] comp1930minVal;
    wire [5:0] comp1930minI, comp1930minJ;
    Comparator comp1930(comp136minVal, comp136minI, comp136minJ, comp137minVal, comp137minI, comp137minJ, comp1930minVal, comp1930minI, comp1930minJ);
    wire [11:0] comp1931minVal;
    wire [5:0] comp1931minI, comp1931minJ;
    Comparator comp1931(comp138minVal, comp138minI, comp138minJ, comp139minVal, comp139minI, comp139minJ, comp1931minVal, comp1931minI, comp1931minJ);
    wire [11:0] comp1932minVal;
    wire [5:0] comp1932minI, comp1932minJ;
    Comparator comp1932(comp140minVal, comp140minI, comp140minJ, comp141minVal, comp141minI, comp141minJ, comp1932minVal, comp1932minI, comp1932minJ);
    wire [11:0] comp1933minVal;
    wire [5:0] comp1933minI, comp1933minJ;
    Comparator comp1933(comp142minVal, comp142minI, comp142minJ, comp143minVal, comp143minI, comp143minJ, comp1933minVal, comp1933minI, comp1933minJ);
    wire [11:0] comp1934minVal;
    wire [5:0] comp1934minI, comp1934minJ;
    Comparator comp1934(comp144minVal, comp144minI, comp144minJ, comp145minVal, comp145minI, comp145minJ, comp1934minVal, comp1934minI, comp1934minJ);
    wire [11:0] comp1935minVal;
    wire [5:0] comp1935minI, comp1935minJ;
    Comparator comp1935(comp146minVal, comp146minI, comp146minJ, comp147minVal, comp147minI, comp147minJ, comp1935minVal, comp1935minI, comp1935minJ);
    wire [11:0] comp1936minVal;
    wire [5:0] comp1936minI, comp1936minJ;
    Comparator comp1936(comp148minVal, comp148minI, comp148minJ, comp149minVal, comp149minI, comp149minJ, comp1936minVal, comp1936minI, comp1936minJ);
    wire [11:0] comp1937minVal;
    wire [5:0] comp1937minI, comp1937minJ;
    Comparator comp1937(comp150minVal, comp150minI, comp150minJ, comp151minVal, comp151minI, comp151minJ, comp1937minVal, comp1937minI, comp1937minJ);
    wire [11:0] comp1938minVal;
    wire [5:0] comp1938minI, comp1938minJ;
    Comparator comp1938(comp152minVal, comp152minI, comp152minJ, comp153minVal, comp153minI, comp153minJ, comp1938minVal, comp1938minI, comp1938minJ);
    wire [11:0] comp1939minVal;
    wire [5:0] comp1939minI, comp1939minJ;
    Comparator comp1939(comp154minVal, comp154minI, comp154minJ, comp155minVal, comp155minI, comp155minJ, comp1939minVal, comp1939minI, comp1939minJ);
    wire [11:0] comp1940minVal;
    wire [5:0] comp1940minI, comp1940minJ;
    Comparator comp1940(comp156minVal, comp156minI, comp156minJ, comp157minVal, comp157minI, comp157minJ, comp1940minVal, comp1940minI, comp1940minJ);
    wire [11:0] comp1941minVal;
    wire [5:0] comp1941minI, comp1941minJ;
    Comparator comp1941(comp158minVal, comp158minI, comp158minJ, comp159minVal, comp159minI, comp159minJ, comp1941minVal, comp1941minI, comp1941minJ);
    wire [11:0] comp1942minVal;
    wire [5:0] comp1942minI, comp1942minJ;
    Comparator comp1942(comp160minVal, comp160minI, comp160minJ, comp161minVal, comp161minI, comp161minJ, comp1942minVal, comp1942minI, comp1942minJ);
    wire [11:0] comp1943minVal;
    wire [5:0] comp1943minI, comp1943minJ;
    Comparator comp1943(comp162minVal, comp162minI, comp162minJ, comp163minVal, comp163minI, comp163minJ, comp1943minVal, comp1943minI, comp1943minJ);
    wire [11:0] comp1944minVal;
    wire [5:0] comp1944minI, comp1944minJ;
    Comparator comp1944(comp164minVal, comp164minI, comp164minJ, comp165minVal, comp165minI, comp165minJ, comp1944minVal, comp1944minI, comp1944minJ);
    wire [11:0] comp1945minVal;
    wire [5:0] comp1945minI, comp1945minJ;
    Comparator comp1945(comp166minVal, comp166minI, comp166minJ, comp167minVal, comp167minI, comp167minJ, comp1945minVal, comp1945minI, comp1945minJ);
    wire [11:0] comp1946minVal;
    wire [5:0] comp1946minI, comp1946minJ;
    Comparator comp1946(comp168minVal, comp168minI, comp168minJ, comp169minVal, comp169minI, comp169minJ, comp1946minVal, comp1946minI, comp1946minJ);
    wire [11:0] comp1947minVal;
    wire [5:0] comp1947minI, comp1947minJ;
    Comparator comp1947(comp170minVal, comp170minI, comp170minJ, comp171minVal, comp171minI, comp171minJ, comp1947minVal, comp1947minI, comp1947minJ);
    wire [11:0] comp1948minVal;
    wire [5:0] comp1948minI, comp1948minJ;
    Comparator comp1948(comp172minVal, comp172minI, comp172minJ, comp173minVal, comp173minI, comp173minJ, comp1948minVal, comp1948minI, comp1948minJ);
    wire [11:0] comp1949minVal;
    wire [5:0] comp1949minI, comp1949minJ;
    Comparator comp1949(comp174minVal, comp174minI, comp174minJ, comp175minVal, comp175minI, comp175minJ, comp1949minVal, comp1949minI, comp1949minJ);
    wire [11:0] comp1950minVal;
    wire [5:0] comp1950minI, comp1950minJ;
    Comparator comp1950(comp176minVal, comp176minI, comp176minJ, comp177minVal, comp177minI, comp177minJ, comp1950minVal, comp1950minI, comp1950minJ);
    wire [11:0] comp1951minVal;
    wire [5:0] comp1951minI, comp1951minJ;
    Comparator comp1951(comp178minVal, comp178minI, comp178minJ, comp179minVal, comp179minI, comp179minJ, comp1951minVal, comp1951minI, comp1951minJ);
    wire [11:0] comp1952minVal;
    wire [5:0] comp1952minI, comp1952minJ;
    Comparator comp1952(comp180minVal, comp180minI, comp180minJ, comp181minVal, comp181minI, comp181minJ, comp1952minVal, comp1952minI, comp1952minJ);
    wire [11:0] comp1953minVal;
    wire [5:0] comp1953minI, comp1953minJ;
    Comparator comp1953(comp182minVal, comp182minI, comp182minJ, comp183minVal, comp183minI, comp183minJ, comp1953minVal, comp1953minI, comp1953minJ);
    wire [11:0] comp1954minVal;
    wire [5:0] comp1954minI, comp1954minJ;
    Comparator comp1954(comp184minVal, comp184minI, comp184minJ, comp185minVal, comp185minI, comp185minJ, comp1954minVal, comp1954minI, comp1954minJ);
    wire [11:0] comp1955minVal;
    wire [5:0] comp1955minI, comp1955minJ;
    Comparator comp1955(comp186minVal, comp186minI, comp186minJ, comp187minVal, comp187minI, comp187minJ, comp1955minVal, comp1955minI, comp1955minJ);
    wire [11:0] comp1956minVal;
    wire [5:0] comp1956minI, comp1956minJ;
    Comparator comp1956(comp188minVal, comp188minI, comp188minJ, comp189minVal, comp189minI, comp189minJ, comp1956minVal, comp1956minI, comp1956minJ);
    wire [11:0] comp1957minVal;
    wire [5:0] comp1957minI, comp1957minJ;
    Comparator comp1957(comp190minVal, comp190minI, comp190minJ, comp191minVal, comp191minI, comp191minJ, comp1957minVal, comp1957minI, comp1957minJ);
    wire [11:0] comp1958minVal;
    wire [5:0] comp1958minI, comp1958minJ;
    Comparator comp1958(comp192minVal, comp192minI, comp192minJ, comp193minVal, comp193minI, comp193minJ, comp1958minVal, comp1958minI, comp1958minJ);
    wire [11:0] comp1959minVal;
    wire [5:0] comp1959minI, comp1959minJ;
    Comparator comp1959(comp194minVal, comp194minI, comp194minJ, comp195minVal, comp195minI, comp195minJ, comp1959minVal, comp1959minI, comp1959minJ);
    wire [11:0] comp1960minVal;
    wire [5:0] comp1960minI, comp1960minJ;
    Comparator comp1960(comp196minVal, comp196minI, comp196minJ, comp197minVal, comp197minI, comp197minJ, comp1960minVal, comp1960minI, comp1960minJ);
    wire [11:0] comp1961minVal;
    wire [5:0] comp1961minI, comp1961minJ;
    Comparator comp1961(comp198minVal, comp198minI, comp198minJ, comp199minVal, comp199minI, comp199minJ, comp1961minVal, comp1961minI, comp1961minJ);
    wire [11:0] comp1962minVal;
    wire [5:0] comp1962minI, comp1962minJ;
    Comparator comp1962(comp200minVal, comp200minI, comp200minJ, comp201minVal, comp201minI, comp201minJ, comp1962minVal, comp1962minI, comp1962minJ);
    wire [11:0] comp1963minVal;
    wire [5:0] comp1963minI, comp1963minJ;
    Comparator comp1963(comp202minVal, comp202minI, comp202minJ, comp203minVal, comp203minI, comp203minJ, comp1963minVal, comp1963minI, comp1963minJ);
    wire [11:0] comp1964minVal;
    wire [5:0] comp1964minI, comp1964minJ;
    Comparator comp1964(comp204minVal, comp204minI, comp204minJ, comp205minVal, comp205minI, comp205minJ, comp1964minVal, comp1964minI, comp1964minJ);
    wire [11:0] comp1965minVal;
    wire [5:0] comp1965minI, comp1965minJ;
    Comparator comp1965(comp206minVal, comp206minI, comp206minJ, comp207minVal, comp207minI, comp207minJ, comp1965minVal, comp1965minI, comp1965minJ);
    wire [11:0] comp1966minVal;
    wire [5:0] comp1966minI, comp1966minJ;
    Comparator comp1966(comp208minVal, comp208minI, comp208minJ, comp209minVal, comp209minI, comp209minJ, comp1966minVal, comp1966minI, comp1966minJ);
    wire [11:0] comp1967minVal;
    wire [5:0] comp1967minI, comp1967minJ;
    Comparator comp1967(comp210minVal, comp210minI, comp210minJ, comp211minVal, comp211minI, comp211minJ, comp1967minVal, comp1967minI, comp1967minJ);
    wire [11:0] comp1968minVal;
    wire [5:0] comp1968minI, comp1968minJ;
    Comparator comp1968(comp212minVal, comp212minI, comp212minJ, comp213minVal, comp213minI, comp213minJ, comp1968minVal, comp1968minI, comp1968minJ);
    wire [11:0] comp1969minVal;
    wire [5:0] comp1969minI, comp1969minJ;
    Comparator comp1969(comp214minVal, comp214minI, comp214minJ, comp215minVal, comp215minI, comp215minJ, comp1969minVal, comp1969minI, comp1969minJ);
    wire [11:0] comp1970minVal;
    wire [5:0] comp1970minI, comp1970minJ;
    Comparator comp1970(comp216minVal, comp216minI, comp216minJ, comp217minVal, comp217minI, comp217minJ, comp1970minVal, comp1970minI, comp1970minJ);
    wire [11:0] comp1971minVal;
    wire [5:0] comp1971minI, comp1971minJ;
    Comparator comp1971(comp218minVal, comp218minI, comp218minJ, comp219minVal, comp219minI, comp219minJ, comp1971minVal, comp1971minI, comp1971minJ);
    wire [11:0] comp1972minVal;
    wire [5:0] comp1972minI, comp1972minJ;
    Comparator comp1972(comp220minVal, comp220minI, comp220minJ, comp221minVal, comp221minI, comp221minJ, comp1972minVal, comp1972minI, comp1972minJ);
    wire [11:0] comp1973minVal;
    wire [5:0] comp1973minI, comp1973minJ;
    Comparator comp1973(comp222minVal, comp222minI, comp222minJ, comp223minVal, comp223minI, comp223minJ, comp1973minVal, comp1973minI, comp1973minJ);
    wire [11:0] comp1974minVal;
    wire [5:0] comp1974minI, comp1974minJ;
    Comparator comp1974(comp224minVal, comp224minI, comp224minJ, comp225minVal, comp225minI, comp225minJ, comp1974minVal, comp1974minI, comp1974minJ);
    wire [11:0] comp1975minVal;
    wire [5:0] comp1975minI, comp1975minJ;
    Comparator comp1975(comp226minVal, comp226minI, comp226minJ, comp227minVal, comp227minI, comp227minJ, comp1975minVal, comp1975minI, comp1975minJ);
    wire [11:0] comp1976minVal;
    wire [5:0] comp1976minI, comp1976minJ;
    Comparator comp1976(comp228minVal, comp228minI, comp228minJ, comp229minVal, comp229minI, comp229minJ, comp1976minVal, comp1976minI, comp1976minJ);
    wire [11:0] comp1977minVal;
    wire [5:0] comp1977minI, comp1977minJ;
    Comparator comp1977(comp230minVal, comp230minI, comp230minJ, comp231minVal, comp231minI, comp231minJ, comp1977minVal, comp1977minI, comp1977minJ);
    wire [11:0] comp1978minVal;
    wire [5:0] comp1978minI, comp1978minJ;
    Comparator comp1978(comp232minVal, comp232minI, comp232minJ, comp233minVal, comp233minI, comp233minJ, comp1978minVal, comp1978minI, comp1978minJ);
    wire [11:0] comp1979minVal;
    wire [5:0] comp1979minI, comp1979minJ;
    Comparator comp1979(comp234minVal, comp234minI, comp234minJ, comp235minVal, comp235minI, comp235minJ, comp1979minVal, comp1979minI, comp1979minJ);
    wire [11:0] comp1980minVal;
    wire [5:0] comp1980minI, comp1980minJ;
    Comparator comp1980(comp236minVal, comp236minI, comp236minJ, comp237minVal, comp237minI, comp237minJ, comp1980minVal, comp1980minI, comp1980minJ);
    wire [11:0] comp1981minVal;
    wire [5:0] comp1981minI, comp1981minJ;
    Comparator comp1981(comp238minVal, comp238minI, comp238minJ, comp239minVal, comp239minI, comp239minJ, comp1981minVal, comp1981minI, comp1981minJ);
    wire [11:0] comp1982minVal;
    wire [5:0] comp1982minI, comp1982minJ;
    Comparator comp1982(comp240minVal, comp240minI, comp240minJ, comp241minVal, comp241minI, comp241minJ, comp1982minVal, comp1982minI, comp1982minJ);
    wire [11:0] comp1983minVal;
    wire [5:0] comp1983minI, comp1983minJ;
    Comparator comp1983(comp242minVal, comp242minI, comp242minJ, comp243minVal, comp243minI, comp243minJ, comp1983minVal, comp1983minI, comp1983minJ);
    wire [11:0] comp1984minVal;
    wire [5:0] comp1984minI, comp1984minJ;
    Comparator comp1984(comp244minVal, comp244minI, comp244minJ, comp245minVal, comp245minI, comp245minJ, comp1984minVal, comp1984minI, comp1984minJ);
    wire [11:0] comp1985minVal;
    wire [5:0] comp1985minI, comp1985minJ;
    Comparator comp1985(comp246minVal, comp246minI, comp246minJ, comp247minVal, comp247minI, comp247minJ, comp1985minVal, comp1985minI, comp1985minJ);
    wire [11:0] comp1986minVal;
    wire [5:0] comp1986minI, comp1986minJ;
    Comparator comp1986(comp248minVal, comp248minI, comp248minJ, comp249minVal, comp249minI, comp249minJ, comp1986minVal, comp1986minI, comp1986minJ);
    wire [11:0] comp1987minVal;
    wire [5:0] comp1987minI, comp1987minJ;
    Comparator comp1987(comp250minVal, comp250minI, comp250minJ, comp251minVal, comp251minI, comp251minJ, comp1987minVal, comp1987minI, comp1987minJ);
    wire [11:0] comp1988minVal;
    wire [5:0] comp1988minI, comp1988minJ;
    Comparator comp1988(comp252minVal, comp252minI, comp252minJ, comp253minVal, comp253minI, comp253minJ, comp1988minVal, comp1988minI, comp1988minJ);
    wire [11:0] comp1989minVal;
    wire [5:0] comp1989minI, comp1989minJ;
    Comparator comp1989(comp254minVal, comp254minI, comp254minJ, comp255minVal, comp255minI, comp255minJ, comp1989minVal, comp1989minI, comp1989minJ);
    wire [11:0] comp1990minVal;
    wire [5:0] comp1990minI, comp1990minJ;
    Comparator comp1990(comp256minVal, comp256minI, comp256minJ, comp257minVal, comp257minI, comp257minJ, comp1990minVal, comp1990minI, comp1990minJ);
    wire [11:0] comp1991minVal;
    wire [5:0] comp1991minI, comp1991minJ;
    Comparator comp1991(comp258minVal, comp258minI, comp258minJ, comp259minVal, comp259minI, comp259minJ, comp1991minVal, comp1991minI, comp1991minJ);
    wire [11:0] comp1992minVal;
    wire [5:0] comp1992minI, comp1992minJ;
    Comparator comp1992(comp260minVal, comp260minI, comp260minJ, comp261minVal, comp261minI, comp261minJ, comp1992minVal, comp1992minI, comp1992minJ);
    wire [11:0] comp1993minVal;
    wire [5:0] comp1993minI, comp1993minJ;
    Comparator comp1993(comp262minVal, comp262minI, comp262minJ, comp263minVal, comp263minI, comp263minJ, comp1993minVal, comp1993minI, comp1993minJ);
    wire [11:0] comp1994minVal;
    wire [5:0] comp1994minI, comp1994minJ;
    Comparator comp1994(comp264minVal, comp264minI, comp264minJ, comp265minVal, comp265minI, comp265minJ, comp1994minVal, comp1994minI, comp1994minJ);
    wire [11:0] comp1995minVal;
    wire [5:0] comp1995minI, comp1995minJ;
    Comparator comp1995(comp266minVal, comp266minI, comp266minJ, comp267minVal, comp267minI, comp267minJ, comp1995minVal, comp1995minI, comp1995minJ);
    wire [11:0] comp1996minVal;
    wire [5:0] comp1996minI, comp1996minJ;
    Comparator comp1996(comp268minVal, comp268minI, comp268minJ, comp269minVal, comp269minI, comp269minJ, comp1996minVal, comp1996minI, comp1996minJ);
    wire [11:0] comp1997minVal;
    wire [5:0] comp1997minI, comp1997minJ;
    Comparator comp1997(comp270minVal, comp270minI, comp270minJ, comp271minVal, comp271minI, comp271minJ, comp1997minVal, comp1997minI, comp1997minJ);
    wire [11:0] comp1998minVal;
    wire [5:0] comp1998minI, comp1998minJ;
    Comparator comp1998(comp272minVal, comp272minI, comp272minJ, comp273minVal, comp273minI, comp273minJ, comp1998minVal, comp1998minI, comp1998minJ);
    wire [11:0] comp1999minVal;
    wire [5:0] comp1999minI, comp1999minJ;
    Comparator comp1999(comp274minVal, comp274minI, comp274minJ, comp275minVal, comp275minI, comp275minJ, comp1999minVal, comp1999minI, comp1999minJ);
    wire [11:0] comp2000minVal;
    wire [5:0] comp2000minI, comp2000minJ;
    Comparator comp2000(comp276minVal, comp276minI, comp276minJ, comp277minVal, comp277minI, comp277minJ, comp2000minVal, comp2000minI, comp2000minJ);
    wire [11:0] comp2001minVal;
    wire [5:0] comp2001minI, comp2001minJ;
    Comparator comp2001(comp278minVal, comp278minI, comp278minJ, comp279minVal, comp279minI, comp279minJ, comp2001minVal, comp2001minI, comp2001minJ);
    wire [11:0] comp2002minVal;
    wire [5:0] comp2002minI, comp2002minJ;
    Comparator comp2002(comp280minVal, comp280minI, comp280minJ, comp281minVal, comp281minI, comp281minJ, comp2002minVal, comp2002minI, comp2002minJ);
    wire [11:0] comp2003minVal;
    wire [5:0] comp2003minI, comp2003minJ;
    Comparator comp2003(comp282minVal, comp282minI, comp282minJ, comp283minVal, comp283minI, comp283minJ, comp2003minVal, comp2003minI, comp2003minJ);
    wire [11:0] comp2004minVal;
    wire [5:0] comp2004minI, comp2004minJ;
    Comparator comp2004(comp284minVal, comp284minI, comp284minJ, comp285minVal, comp285minI, comp285minJ, comp2004minVal, comp2004minI, comp2004minJ);
    wire [11:0] comp2005minVal;
    wire [5:0] comp2005minI, comp2005minJ;
    Comparator comp2005(comp286minVal, comp286minI, comp286minJ, comp287minVal, comp287minI, comp287minJ, comp2005minVal, comp2005minI, comp2005minJ);
    wire [11:0] comp2006minVal;
    wire [5:0] comp2006minI, comp2006minJ;
    Comparator comp2006(comp288minVal, comp288minI, comp288minJ, comp289minVal, comp289minI, comp289minJ, comp2006minVal, comp2006minI, comp2006minJ);
    wire [11:0] comp2007minVal;
    wire [5:0] comp2007minI, comp2007minJ;
    Comparator comp2007(comp290minVal, comp290minI, comp290minJ, comp291minVal, comp291minI, comp291minJ, comp2007minVal, comp2007minI, comp2007minJ);
    wire [11:0] comp2008minVal;
    wire [5:0] comp2008minI, comp2008minJ;
    Comparator comp2008(comp292minVal, comp292minI, comp292minJ, comp293minVal, comp293minI, comp293minJ, comp2008minVal, comp2008minI, comp2008minJ);
    wire [11:0] comp2009minVal;
    wire [5:0] comp2009minI, comp2009minJ;
    Comparator comp2009(comp294minVal, comp294minI, comp294minJ, comp295minVal, comp295minI, comp295minJ, comp2009minVal, comp2009minI, comp2009minJ);
    wire [11:0] comp2010minVal;
    wire [5:0] comp2010minI, comp2010minJ;
    Comparator comp2010(comp296minVal, comp296minI, comp296minJ, comp297minVal, comp297minI, comp297minJ, comp2010minVal, comp2010minI, comp2010minJ);
    wire [11:0] comp2011minVal;
    wire [5:0] comp2011minI, comp2011minJ;
    Comparator comp2011(comp298minVal, comp298minI, comp298minJ, comp299minVal, comp299minI, comp299minJ, comp2011minVal, comp2011minI, comp2011minJ);
    wire [11:0] comp2012minVal;
    wire [5:0] comp2012minI, comp2012minJ;
    Comparator comp2012(comp300minVal, comp300minI, comp300minJ, comp301minVal, comp301minI, comp301minJ, comp2012minVal, comp2012minI, comp2012minJ);
    wire [11:0] comp2013minVal;
    wire [5:0] comp2013minI, comp2013minJ;
    Comparator comp2013(comp302minVal, comp302minI, comp302minJ, comp303minVal, comp303minI, comp303minJ, comp2013minVal, comp2013minI, comp2013minJ);
    wire [11:0] comp2014minVal;
    wire [5:0] comp2014minI, comp2014minJ;
    Comparator comp2014(comp304minVal, comp304minI, comp304minJ, comp305minVal, comp305minI, comp305minJ, comp2014minVal, comp2014minI, comp2014minJ);
    wire [11:0] comp2015minVal;
    wire [5:0] comp2015minI, comp2015minJ;
    Comparator comp2015(comp306minVal, comp306minI, comp306minJ, comp307minVal, comp307minI, comp307minJ, comp2015minVal, comp2015minI, comp2015minJ);
    wire [11:0] comp2016minVal;
    wire [5:0] comp2016minI, comp2016minJ;
    Comparator comp2016(comp308minVal, comp308minI, comp308minJ, comp309minVal, comp309minI, comp309minJ, comp2016minVal, comp2016minI, comp2016minJ);
    wire [11:0] comp2017minVal;
    wire [5:0] comp2017minI, comp2017minJ;
    Comparator comp2017(comp310minVal, comp310minI, comp310minJ, comp311minVal, comp311minI, comp311minJ, comp2017minVal, comp2017minI, comp2017minJ);
    wire [11:0] comp2018minVal;
    wire [5:0] comp2018minI, comp2018minJ;
    Comparator comp2018(comp312minVal, comp312minI, comp312minJ, comp313minVal, comp313minI, comp313minJ, comp2018minVal, comp2018minI, comp2018minJ);
    wire [11:0] comp2019minVal;
    wire [5:0] comp2019minI, comp2019minJ;
    Comparator comp2019(comp314minVal, comp314minI, comp314minJ, comp315minVal, comp315minI, comp315minJ, comp2019minVal, comp2019minI, comp2019minJ);
    wire [11:0] comp2020minVal;
    wire [5:0] comp2020minI, comp2020minJ;
    Comparator comp2020(comp316minVal, comp316minI, comp316minJ, comp317minVal, comp317minI, comp317minJ, comp2020minVal, comp2020minI, comp2020minJ);
    wire [11:0] comp2021minVal;
    wire [5:0] comp2021minI, comp2021minJ;
    Comparator comp2021(comp318minVal, comp318minI, comp318minJ, comp319minVal, comp319minI, comp319minJ, comp2021minVal, comp2021minI, comp2021minJ);
    wire [11:0] comp2022minVal;
    wire [5:0] comp2022minI, comp2022minJ;
    Comparator comp2022(comp320minVal, comp320minI, comp320minJ, comp321minVal, comp321minI, comp321minJ, comp2022minVal, comp2022minI, comp2022minJ);
    wire [11:0] comp2023minVal;
    wire [5:0] comp2023minI, comp2023minJ;
    Comparator comp2023(comp322minVal, comp322minI, comp322minJ, comp323minVal, comp323minI, comp323minJ, comp2023minVal, comp2023minI, comp2023minJ);
    wire [11:0] comp2024minVal;
    wire [5:0] comp2024minI, comp2024minJ;
    Comparator comp2024(comp324minVal, comp324minI, comp324minJ, comp325minVal, comp325minI, comp325minJ, comp2024minVal, comp2024minI, comp2024minJ);
    wire [11:0] comp2025minVal;
    wire [5:0] comp2025minI, comp2025minJ;
    Comparator comp2025(comp326minVal, comp326minI, comp326minJ, comp327minVal, comp327minI, comp327minJ, comp2025minVal, comp2025minI, comp2025minJ);
    wire [11:0] comp2026minVal;
    wire [5:0] comp2026minI, comp2026minJ;
    Comparator comp2026(comp328minVal, comp328minI, comp328minJ, comp329minVal, comp329minI, comp329minJ, comp2026minVal, comp2026minI, comp2026minJ);
    wire [11:0] comp2027minVal;
    wire [5:0] comp2027minI, comp2027minJ;
    Comparator comp2027(comp330minVal, comp330minI, comp330minJ, comp331minVal, comp331minI, comp331minJ, comp2027minVal, comp2027minI, comp2027minJ);
    wire [11:0] comp2028minVal;
    wire [5:0] comp2028minI, comp2028minJ;
    Comparator comp2028(comp332minVal, comp332minI, comp332minJ, comp333minVal, comp333minI, comp333minJ, comp2028minVal, comp2028minI, comp2028minJ);
    wire [11:0] comp2029minVal;
    wire [5:0] comp2029minI, comp2029minJ;
    Comparator comp2029(comp334minVal, comp334minI, comp334minJ, comp335minVal, comp335minI, comp335minJ, comp2029minVal, comp2029minI, comp2029minJ);
    wire [11:0] comp2030minVal;
    wire [5:0] comp2030minI, comp2030minJ;
    Comparator comp2030(comp336minVal, comp336minI, comp336minJ, comp337minVal, comp337minI, comp337minJ, comp2030minVal, comp2030minI, comp2030minJ);
    wire [11:0] comp2031minVal;
    wire [5:0] comp2031minI, comp2031minJ;
    Comparator comp2031(comp338minVal, comp338minI, comp338minJ, comp339minVal, comp339minI, comp339minJ, comp2031minVal, comp2031minI, comp2031minJ);
    wire [11:0] comp2032minVal;
    wire [5:0] comp2032minI, comp2032minJ;
    Comparator comp2032(comp340minVal, comp340minI, comp340minJ, comp341minVal, comp341minI, comp341minJ, comp2032minVal, comp2032minI, comp2032minJ);
    wire [11:0] comp2033minVal;
    wire [5:0] comp2033minI, comp2033minJ;
    Comparator comp2033(comp342minVal, comp342minI, comp342minJ, comp343minVal, comp343minI, comp343minJ, comp2033minVal, comp2033minI, comp2033minJ);
    wire [11:0] comp2034minVal;
    wire [5:0] comp2034minI, comp2034minJ;
    Comparator comp2034(comp344minVal, comp344minI, comp344minJ, comp345minVal, comp345minI, comp345minJ, comp2034minVal, comp2034minI, comp2034minJ);
    wire [11:0] comp2035minVal;
    wire [5:0] comp2035minI, comp2035minJ;
    Comparator comp2035(comp346minVal, comp346minI, comp346minJ, comp347minVal, comp347minI, comp347minJ, comp2035minVal, comp2035minI, comp2035minJ);
    wire [11:0] comp2036minVal;
    wire [5:0] comp2036minI, comp2036minJ;
    Comparator comp2036(comp348minVal, comp348minI, comp348minJ, comp349minVal, comp349minI, comp349minJ, comp2036minVal, comp2036minI, comp2036minJ);
    wire [11:0] comp2037minVal;
    wire [5:0] comp2037minI, comp2037minJ;
    Comparator comp2037(comp350minVal, comp350minI, comp350minJ, comp351minVal, comp351minI, comp351minJ, comp2037minVal, comp2037minI, comp2037minJ);
    wire [11:0] comp2038minVal;
    wire [5:0] comp2038minI, comp2038minJ;
    Comparator comp2038(comp352minVal, comp352minI, comp352minJ, comp353minVal, comp353minI, comp353minJ, comp2038minVal, comp2038minI, comp2038minJ);
    wire [11:0] comp2039minVal;
    wire [5:0] comp2039minI, comp2039minJ;
    Comparator comp2039(comp354minVal, comp354minI, comp354minJ, comp355minVal, comp355minI, comp355minJ, comp2039minVal, comp2039minI, comp2039minJ);
    wire [11:0] comp2040minVal;
    wire [5:0] comp2040minI, comp2040minJ;
    Comparator comp2040(comp356minVal, comp356minI, comp356minJ, comp357minVal, comp357minI, comp357minJ, comp2040minVal, comp2040minI, comp2040minJ);
    wire [11:0] comp2041minVal;
    wire [5:0] comp2041minI, comp2041minJ;
    Comparator comp2041(comp358minVal, comp358minI, comp358minJ, comp359minVal, comp359minI, comp359minJ, comp2041minVal, comp2041minI, comp2041minJ);
    wire [11:0] comp2042minVal;
    wire [5:0] comp2042minI, comp2042minJ;
    Comparator comp2042(comp360minVal, comp360minI, comp360minJ, comp361minVal, comp361minI, comp361minJ, comp2042minVal, comp2042minI, comp2042minJ);
    wire [11:0] comp2043minVal;
    wire [5:0] comp2043minI, comp2043minJ;
    Comparator comp2043(comp362minVal, comp362minI, comp362minJ, comp363minVal, comp363minI, comp363minJ, comp2043minVal, comp2043minI, comp2043minJ);
    wire [11:0] comp2044minVal;
    wire [5:0] comp2044minI, comp2044minJ;
    Comparator comp2044(comp364minVal, comp364minI, comp364minJ, comp365minVal, comp365minI, comp365minJ, comp2044minVal, comp2044minI, comp2044minJ);
    wire [11:0] comp2045minVal;
    wire [5:0] comp2045minI, comp2045minJ;
    Comparator comp2045(comp366minVal, comp366minI, comp366minJ, comp367minVal, comp367minI, comp367minJ, comp2045minVal, comp2045minI, comp2045minJ);
    wire [11:0] comp2046minVal;
    wire [5:0] comp2046minI, comp2046minJ;
    Comparator comp2046(comp368minVal, comp368minI, comp368minJ, comp369minVal, comp369minI, comp369minJ, comp2046minVal, comp2046minI, comp2046minJ);
    wire [11:0] comp2047minVal;
    wire [5:0] comp2047minI, comp2047minJ;
    Comparator comp2047(comp370minVal, comp370minI, comp370minJ, comp371minVal, comp371minI, comp371minJ, comp2047minVal, comp2047minI, comp2047minJ);
    wire [11:0] comp2048minVal;
    wire [5:0] comp2048minI, comp2048minJ;
    Comparator comp2048(comp372minVal, comp372minI, comp372minJ, comp373minVal, comp373minI, comp373minJ, comp2048minVal, comp2048minI, comp2048minJ);
    wire [11:0] comp2049minVal;
    wire [5:0] comp2049minI, comp2049minJ;
    Comparator comp2049(comp374minVal, comp374minI, comp374minJ, comp375minVal, comp375minI, comp375minJ, comp2049minVal, comp2049minI, comp2049minJ);
    wire [11:0] comp2050minVal;
    wire [5:0] comp2050minI, comp2050minJ;
    Comparator comp2050(comp376minVal, comp376minI, comp376minJ, comp377minVal, comp377minI, comp377minJ, comp2050minVal, comp2050minI, comp2050minJ);
    wire [11:0] comp2051minVal;
    wire [5:0] comp2051minI, comp2051minJ;
    Comparator comp2051(comp378minVal, comp378minI, comp378minJ, comp379minVal, comp379minI, comp379minJ, comp2051minVal, comp2051minI, comp2051minJ);
    wire [11:0] comp2052minVal;
    wire [5:0] comp2052minI, comp2052minJ;
    Comparator comp2052(comp380minVal, comp380minI, comp380minJ, comp381minVal, comp381minI, comp381minJ, comp2052minVal, comp2052minI, comp2052minJ);
    wire [11:0] comp2053minVal;
    wire [5:0] comp2053minI, comp2053minJ;
    Comparator comp2053(comp382minVal, comp382minI, comp382minJ, comp383minVal, comp383minI, comp383minJ, comp2053minVal, comp2053minI, comp2053minJ);
    wire [11:0] comp2054minVal;
    wire [5:0] comp2054minI, comp2054minJ;
    Comparator comp2054(comp384minVal, comp384minI, comp384minJ, comp385minVal, comp385minI, comp385minJ, comp2054minVal, comp2054minI, comp2054minJ);
    wire [11:0] comp2055minVal;
    wire [5:0] comp2055minI, comp2055minJ;
    Comparator comp2055(comp386minVal, comp386minI, comp386minJ, comp387minVal, comp387minI, comp387minJ, comp2055minVal, comp2055minI, comp2055minJ);
    wire [11:0] comp2056minVal;
    wire [5:0] comp2056minI, comp2056minJ;
    Comparator comp2056(comp388minVal, comp388minI, comp388minJ, comp389minVal, comp389minI, comp389minJ, comp2056minVal, comp2056minI, comp2056minJ);
    wire [11:0] comp2057minVal;
    wire [5:0] comp2057minI, comp2057minJ;
    Comparator comp2057(comp390minVal, comp390minI, comp390minJ, comp391minVal, comp391minI, comp391minJ, comp2057minVal, comp2057minI, comp2057minJ);
    wire [11:0] comp2058minVal;
    wire [5:0] comp2058minI, comp2058minJ;
    Comparator comp2058(comp392minVal, comp392minI, comp392minJ, comp393minVal, comp393minI, comp393minJ, comp2058minVal, comp2058minI, comp2058minJ);
    wire [11:0] comp2059minVal;
    wire [5:0] comp2059minI, comp2059minJ;
    Comparator comp2059(comp394minVal, comp394minI, comp394minJ, comp395minVal, comp395minI, comp395minJ, comp2059minVal, comp2059minI, comp2059minJ);
    wire [11:0] comp2060minVal;
    wire [5:0] comp2060minI, comp2060minJ;
    Comparator comp2060(comp396minVal, comp396minI, comp396minJ, comp397minVal, comp397minI, comp397minJ, comp2060minVal, comp2060minI, comp2060minJ);
    wire [11:0] comp2061minVal;
    wire [5:0] comp2061minI, comp2061minJ;
    Comparator comp2061(comp398minVal, comp398minI, comp398minJ, comp399minVal, comp399minI, comp399minJ, comp2061minVal, comp2061minI, comp2061minJ);
    wire [11:0] comp2062minVal;
    wire [5:0] comp2062minI, comp2062minJ;
    Comparator comp2062(comp400minVal, comp400minI, comp400minJ, comp401minVal, comp401minI, comp401minJ, comp2062minVal, comp2062minI, comp2062minJ);
    wire [11:0] comp2063minVal;
    wire [5:0] comp2063minI, comp2063minJ;
    Comparator comp2063(comp402minVal, comp402minI, comp402minJ, comp403minVal, comp403minI, comp403minJ, comp2063minVal, comp2063minI, comp2063minJ);
    wire [11:0] comp2064minVal;
    wire [5:0] comp2064minI, comp2064minJ;
    Comparator comp2064(comp404minVal, comp404minI, comp404minJ, comp405minVal, comp405minI, comp405minJ, comp2064minVal, comp2064minI, comp2064minJ);
    wire [11:0] comp2065minVal;
    wire [5:0] comp2065minI, comp2065minJ;
    Comparator comp2065(comp406minVal, comp406minI, comp406minJ, comp407minVal, comp407minI, comp407minJ, comp2065minVal, comp2065minI, comp2065minJ);
    wire [11:0] comp2066minVal;
    wire [5:0] comp2066minI, comp2066minJ;
    Comparator comp2066(comp408minVal, comp408minI, comp408minJ, comp409minVal, comp409minI, comp409minJ, comp2066minVal, comp2066minI, comp2066minJ);
    wire [11:0] comp2067minVal;
    wire [5:0] comp2067minI, comp2067minJ;
    Comparator comp2067(comp410minVal, comp410minI, comp410minJ, comp411minVal, comp411minI, comp411minJ, comp2067minVal, comp2067minI, comp2067minJ);
    wire [11:0] comp2068minVal;
    wire [5:0] comp2068minI, comp2068minJ;
    Comparator comp2068(comp412minVal, comp412minI, comp412minJ, comp413minVal, comp413minI, comp413minJ, comp2068minVal, comp2068minI, comp2068minJ);
    wire [11:0] comp2069minVal;
    wire [5:0] comp2069minI, comp2069minJ;
    Comparator comp2069(comp414minVal, comp414minI, comp414minJ, comp415minVal, comp415minI, comp415minJ, comp2069minVal, comp2069minI, comp2069minJ);
    wire [11:0] comp2070minVal;
    wire [5:0] comp2070minI, comp2070minJ;
    Comparator comp2070(comp416minVal, comp416minI, comp416minJ, comp417minVal, comp417minI, comp417minJ, comp2070minVal, comp2070minI, comp2070minJ);
    wire [11:0] comp2071minVal;
    wire [5:0] comp2071minI, comp2071minJ;
    Comparator comp2071(comp418minVal, comp418minI, comp418minJ, comp419minVal, comp419minI, comp419minJ, comp2071minVal, comp2071minI, comp2071minJ);
    wire [11:0] comp2072minVal;
    wire [5:0] comp2072minI, comp2072minJ;
    Comparator comp2072(comp420minVal, comp420minI, comp420minJ, comp421minVal, comp421minI, comp421minJ, comp2072minVal, comp2072minI, comp2072minJ);
    wire [11:0] comp2073minVal;
    wire [5:0] comp2073minI, comp2073minJ;
    Comparator comp2073(comp422minVal, comp422minI, comp422minJ, comp423minVal, comp423minI, comp423minJ, comp2073minVal, comp2073minI, comp2073minJ);
    wire [11:0] comp2074minVal;
    wire [5:0] comp2074minI, comp2074minJ;
    Comparator comp2074(comp424minVal, comp424minI, comp424minJ, comp425minVal, comp425minI, comp425minJ, comp2074minVal, comp2074minI, comp2074minJ);
    wire [11:0] comp2075minVal;
    wire [5:0] comp2075minI, comp2075minJ;
    Comparator comp2075(comp426minVal, comp426minI, comp426minJ, comp427minVal, comp427minI, comp427minJ, comp2075minVal, comp2075minI, comp2075minJ);
    wire [11:0] comp2076minVal;
    wire [5:0] comp2076minI, comp2076minJ;
    Comparator comp2076(comp428minVal, comp428minI, comp428minJ, comp429minVal, comp429minI, comp429minJ, comp2076minVal, comp2076minI, comp2076minJ);
    wire [11:0] comp2077minVal;
    wire [5:0] comp2077minI, comp2077minJ;
    Comparator comp2077(comp430minVal, comp430minI, comp430minJ, comp431minVal, comp431minI, comp431minJ, comp2077minVal, comp2077minI, comp2077minJ);
    wire [11:0] comp2078minVal;
    wire [5:0] comp2078minI, comp2078minJ;
    Comparator comp2078(comp432minVal, comp432minI, comp432minJ, comp433minVal, comp433minI, comp433minJ, comp2078minVal, comp2078minI, comp2078minJ);
    wire [11:0] comp2079minVal;
    wire [5:0] comp2079minI, comp2079minJ;
    Comparator comp2079(comp434minVal, comp434minI, comp434minJ, comp435minVal, comp435minI, comp435minJ, comp2079minVal, comp2079minI, comp2079minJ);
    wire [11:0] comp2080minVal;
    wire [5:0] comp2080minI, comp2080minJ;
    Comparator comp2080(comp436minVal, comp436minI, comp436minJ, comp437minVal, comp437minI, comp437minJ, comp2080minVal, comp2080minI, comp2080minJ);
    wire [11:0] comp2081minVal;
    wire [5:0] comp2081minI, comp2081minJ;
    Comparator comp2081(comp438minVal, comp438minI, comp438minJ, comp439minVal, comp439minI, comp439minJ, comp2081minVal, comp2081minI, comp2081minJ);
    wire [11:0] comp2082minVal;
    wire [5:0] comp2082minI, comp2082minJ;
    Comparator comp2082(comp440minVal, comp440minI, comp440minJ, comp441minVal, comp441minI, comp441minJ, comp2082minVal, comp2082minI, comp2082minJ);
    wire [11:0] comp2083minVal;
    wire [5:0] comp2083minI, comp2083minJ;
    Comparator comp2083(comp442minVal, comp442minI, comp442minJ, comp443minVal, comp443minI, comp443minJ, comp2083minVal, comp2083minI, comp2083minJ);
    wire [11:0] comp2084minVal;
    wire [5:0] comp2084minI, comp2084minJ;
    Comparator comp2084(comp444minVal, comp444minI, comp444minJ, comp445minVal, comp445minI, comp445minJ, comp2084minVal, comp2084minI, comp2084minJ);
    wire [11:0] comp2085minVal;
    wire [5:0] comp2085minI, comp2085minJ;
    Comparator comp2085(comp446minVal, comp446minI, comp446minJ, comp447minVal, comp447minI, comp447minJ, comp2085minVal, comp2085minI, comp2085minJ);
    wire [11:0] comp2086minVal;
    wire [5:0] comp2086minI, comp2086minJ;
    Comparator comp2086(comp448minVal, comp448minI, comp448minJ, comp449minVal, comp449minI, comp449minJ, comp2086minVal, comp2086minI, comp2086minJ);
    wire [11:0] comp2087minVal;
    wire [5:0] comp2087minI, comp2087minJ;
    Comparator comp2087(comp450minVal, comp450minI, comp450minJ, comp451minVal, comp451minI, comp451minJ, comp2087minVal, comp2087minI, comp2087minJ);
    wire [11:0] comp2088minVal;
    wire [5:0] comp2088minI, comp2088minJ;
    Comparator comp2088(comp452minVal, comp452minI, comp452minJ, comp453minVal, comp453minI, comp453minJ, comp2088minVal, comp2088minI, comp2088minJ);
    wire [11:0] comp2089minVal;
    wire [5:0] comp2089minI, comp2089minJ;
    Comparator comp2089(comp454minVal, comp454minI, comp454minJ, comp455minVal, comp455minI, comp455minJ, comp2089minVal, comp2089minI, comp2089minJ);
    wire [11:0] comp2090minVal;
    wire [5:0] comp2090minI, comp2090minJ;
    Comparator comp2090(comp456minVal, comp456minI, comp456minJ, comp457minVal, comp457minI, comp457minJ, comp2090minVal, comp2090minI, comp2090minJ);
    wire [11:0] comp2091minVal;
    wire [5:0] comp2091minI, comp2091minJ;
    Comparator comp2091(comp458minVal, comp458minI, comp458minJ, comp459minVal, comp459minI, comp459minJ, comp2091minVal, comp2091minI, comp2091minJ);
    wire [11:0] comp2092minVal;
    wire [5:0] comp2092minI, comp2092minJ;
    Comparator comp2092(comp460minVal, comp460minI, comp460minJ, comp461minVal, comp461minI, comp461minJ, comp2092minVal, comp2092minI, comp2092minJ);
    wire [11:0] comp2093minVal;
    wire [5:0] comp2093minI, comp2093minJ;
    Comparator comp2093(comp462minVal, comp462minI, comp462minJ, comp463minVal, comp463minI, comp463minJ, comp2093minVal, comp2093minI, comp2093minJ);
    wire [11:0] comp2094minVal;
    wire [5:0] comp2094minI, comp2094minJ;
    Comparator comp2094(comp464minVal, comp464minI, comp464minJ, comp465minVal, comp465minI, comp465minJ, comp2094minVal, comp2094minI, comp2094minJ);
    wire [11:0] comp2095minVal;
    wire [5:0] comp2095minI, comp2095minJ;
    Comparator comp2095(comp466minVal, comp466minI, comp466minJ, comp467minVal, comp467minI, comp467minJ, comp2095minVal, comp2095minI, comp2095minJ);
    wire [11:0] comp2096minVal;
    wire [5:0] comp2096minI, comp2096minJ;
    Comparator comp2096(comp468minVal, comp468minI, comp468minJ, comp469minVal, comp469minI, comp469minJ, comp2096minVal, comp2096minI, comp2096minJ);
    wire [11:0] comp2097minVal;
    wire [5:0] comp2097minI, comp2097minJ;
    Comparator comp2097(comp470minVal, comp470minI, comp470minJ, comp471minVal, comp471minI, comp471minJ, comp2097minVal, comp2097minI, comp2097minJ);
    wire [11:0] comp2098minVal;
    wire [5:0] comp2098minI, comp2098minJ;
    Comparator comp2098(comp472minVal, comp472minI, comp472minJ, comp473minVal, comp473minI, comp473minJ, comp2098minVal, comp2098minI, comp2098minJ);
    wire [11:0] comp2099minVal;
    wire [5:0] comp2099minI, comp2099minJ;
    Comparator comp2099(comp474minVal, comp474minI, comp474minJ, comp475minVal, comp475minI, comp475minJ, comp2099minVal, comp2099minI, comp2099minJ);
    wire [11:0] comp2100minVal;
    wire [5:0] comp2100minI, comp2100minJ;
    Comparator comp2100(comp476minVal, comp476minI, comp476minJ, comp477minVal, comp477minI, comp477minJ, comp2100minVal, comp2100minI, comp2100minJ);
    wire [11:0] comp2101minVal;
    wire [5:0] comp2101minI, comp2101minJ;
    Comparator comp2101(comp478minVal, comp478minI, comp478minJ, comp479minVal, comp479minI, comp479minJ, comp2101minVal, comp2101minI, comp2101minJ);
    wire [11:0] comp2102minVal;
    wire [5:0] comp2102minI, comp2102minJ;
    Comparator comp2102(comp480minVal, comp480minI, comp480minJ, comp481minVal, comp481minI, comp481minJ, comp2102minVal, comp2102minI, comp2102minJ);
    wire [11:0] comp2103minVal;
    wire [5:0] comp2103minI, comp2103minJ;
    Comparator comp2103(comp482minVal, comp482minI, comp482minJ, comp483minVal, comp483minI, comp483minJ, comp2103minVal, comp2103minI, comp2103minJ);
    wire [11:0] comp2104minVal;
    wire [5:0] comp2104minI, comp2104minJ;
    Comparator comp2104(comp484minVal, comp484minI, comp484minJ, comp485minVal, comp485minI, comp485minJ, comp2104minVal, comp2104minI, comp2104minJ);
    wire [11:0] comp2105minVal;
    wire [5:0] comp2105minI, comp2105minJ;
    Comparator comp2105(comp486minVal, comp486minI, comp486minJ, comp487minVal, comp487minI, comp487minJ, comp2105minVal, comp2105minI, comp2105minJ);
    wire [11:0] comp2106minVal;
    wire [5:0] comp2106minI, comp2106minJ;
    Comparator comp2106(comp488minVal, comp488minI, comp488minJ, comp489minVal, comp489minI, comp489minJ, comp2106minVal, comp2106minI, comp2106minJ);
    wire [11:0] comp2107minVal;
    wire [5:0] comp2107minI, comp2107minJ;
    Comparator comp2107(comp490minVal, comp490minI, comp490minJ, comp491minVal, comp491minI, comp491minJ, comp2107minVal, comp2107minI, comp2107minJ);
    wire [11:0] comp2108minVal;
    wire [5:0] comp2108minI, comp2108minJ;
    Comparator comp2108(comp492minVal, comp492minI, comp492minJ, comp493minVal, comp493minI, comp493minJ, comp2108minVal, comp2108minI, comp2108minJ);
    wire [11:0] comp2109minVal;
    wire [5:0] comp2109minI, comp2109minJ;
    Comparator comp2109(comp494minVal, comp494minI, comp494minJ, comp495minVal, comp495minI, comp495minJ, comp2109minVal, comp2109minI, comp2109minJ);
    wire [11:0] comp2110minVal;
    wire [5:0] comp2110minI, comp2110minJ;
    Comparator comp2110(comp496minVal, comp496minI, comp496minJ, comp497minVal, comp497minI, comp497minJ, comp2110minVal, comp2110minI, comp2110minJ);
    wire [11:0] comp2111minVal;
    wire [5:0] comp2111minI, comp2111minJ;
    Comparator comp2111(comp498minVal, comp498minI, comp498minJ, comp499minVal, comp499minI, comp499minJ, comp2111minVal, comp2111minI, comp2111minJ);
    wire [11:0] comp2112minVal;
    wire [5:0] comp2112minI, comp2112minJ;
    Comparator comp2112(comp500minVal, comp500minI, comp500minJ, comp501minVal, comp501minI, comp501minJ, comp2112minVal, comp2112minI, comp2112minJ);
    wire [11:0] comp2113minVal;
    wire [5:0] comp2113minI, comp2113minJ;
    Comparator comp2113(comp502minVal, comp502minI, comp502minJ, comp503minVal, comp503minI, comp503minJ, comp2113minVal, comp2113minI, comp2113minJ);
    wire [11:0] comp2114minVal;
    wire [5:0] comp2114minI, comp2114minJ;
    Comparator comp2114(comp504minVal, comp504minI, comp504minJ, comp505minVal, comp505minI, comp505minJ, comp2114minVal, comp2114minI, comp2114minJ);
    wire [11:0] comp2115minVal;
    wire [5:0] comp2115minI, comp2115minJ;
    Comparator comp2115(comp506minVal, comp506minI, comp506minJ, comp507minVal, comp507minI, comp507minJ, comp2115minVal, comp2115minI, comp2115minJ);
    wire [11:0] comp2116minVal;
    wire [5:0] comp2116minI, comp2116minJ;
    Comparator comp2116(comp508minVal, comp508minI, comp508minJ, comp509minVal, comp509minI, comp509minJ, comp2116minVal, comp2116minI, comp2116minJ);
    wire [11:0] comp2117minVal;
    wire [5:0] comp2117minI, comp2117minJ;
    Comparator comp2117(comp510minVal, comp510minI, comp510minJ, comp511minVal, comp511minI, comp511minJ, comp2117minVal, comp2117minI, comp2117minJ);
    wire [11:0] comp2118minVal;
    wire [5:0] comp2118minI, comp2118minJ;
    Comparator comp2118(comp512minVal, comp512minI, comp512minJ, comp513minVal, comp513minI, comp513minJ, comp2118minVal, comp2118minI, comp2118minJ);
    wire [11:0] comp2119minVal;
    wire [5:0] comp2119minI, comp2119minJ;
    Comparator comp2119(comp514minVal, comp514minI, comp514minJ, comp515minVal, comp515minI, comp515minJ, comp2119minVal, comp2119minI, comp2119minJ);
    wire [11:0] comp2120minVal;
    wire [5:0] comp2120minI, comp2120minJ;
    Comparator comp2120(comp516minVal, comp516minI, comp516minJ, comp517minVal, comp517minI, comp517minJ, comp2120minVal, comp2120minI, comp2120minJ);
    wire [11:0] comp2121minVal;
    wire [5:0] comp2121minI, comp2121minJ;
    Comparator comp2121(comp518minVal, comp518minI, comp518minJ, comp519minVal, comp519minI, comp519minJ, comp2121minVal, comp2121minI, comp2121minJ);
    wire [11:0] comp2122minVal;
    wire [5:0] comp2122minI, comp2122minJ;
    Comparator comp2122(comp520minVal, comp520minI, comp520minJ, comp521minVal, comp521minI, comp521minJ, comp2122minVal, comp2122minI, comp2122minJ);
    wire [11:0] comp2123minVal;
    wire [5:0] comp2123minI, comp2123minJ;
    Comparator comp2123(comp522minVal, comp522minI, comp522minJ, comp523minVal, comp523minI, comp523minJ, comp2123minVal, comp2123minI, comp2123minJ);
    wire [11:0] comp2124minVal;
    wire [5:0] comp2124minI, comp2124minJ;
    Comparator comp2124(comp524minVal, comp524minI, comp524minJ, comp525minVal, comp525minI, comp525minJ, comp2124minVal, comp2124minI, comp2124minJ);
    wire [11:0] comp2125minVal;
    wire [5:0] comp2125minI, comp2125minJ;
    Comparator comp2125(comp526minVal, comp526minI, comp526minJ, comp527minVal, comp527minI, comp527minJ, comp2125minVal, comp2125minI, comp2125minJ);
    wire [11:0] comp2126minVal;
    wire [5:0] comp2126minI, comp2126minJ;
    Comparator comp2126(comp528minVal, comp528minI, comp528minJ, comp529minVal, comp529minI, comp529minJ, comp2126minVal, comp2126minI, comp2126minJ);
    wire [11:0] comp2127minVal;
    wire [5:0] comp2127minI, comp2127minJ;
    Comparator comp2127(comp530minVal, comp530minI, comp530minJ, comp531minVal, comp531minI, comp531minJ, comp2127minVal, comp2127minI, comp2127minJ);
    wire [11:0] comp2128minVal;
    wire [5:0] comp2128minI, comp2128minJ;
    Comparator comp2128(comp532minVal, comp532minI, comp532minJ, comp533minVal, comp533minI, comp533minJ, comp2128minVal, comp2128minI, comp2128minJ);
    wire [11:0] comp2129minVal;
    wire [5:0] comp2129minI, comp2129minJ;
    Comparator comp2129(comp534minVal, comp534minI, comp534minJ, comp535minVal, comp535minI, comp535minJ, comp2129minVal, comp2129minI, comp2129minJ);
    wire [11:0] comp2130minVal;
    wire [5:0] comp2130minI, comp2130minJ;
    Comparator comp2130(comp536minVal, comp536minI, comp536minJ, comp537minVal, comp537minI, comp537minJ, comp2130minVal, comp2130minI, comp2130minJ);
    wire [11:0] comp2131minVal;
    wire [5:0] comp2131minI, comp2131minJ;
    Comparator comp2131(comp538minVal, comp538minI, comp538minJ, comp539minVal, comp539minI, comp539minJ, comp2131minVal, comp2131minI, comp2131minJ);
    wire [11:0] comp2132minVal;
    wire [5:0] comp2132minI, comp2132minJ;
    Comparator comp2132(comp540minVal, comp540minI, comp540minJ, comp541minVal, comp541minI, comp541minJ, comp2132minVal, comp2132minI, comp2132minJ);
    wire [11:0] comp2133minVal;
    wire [5:0] comp2133minI, comp2133minJ;
    Comparator comp2133(comp542minVal, comp542minI, comp542minJ, comp543minVal, comp543minI, comp543minJ, comp2133minVal, comp2133minI, comp2133minJ);
    wire [11:0] comp2134minVal;
    wire [5:0] comp2134minI, comp2134minJ;
    Comparator comp2134(comp544minVal, comp544minI, comp544minJ, comp545minVal, comp545minI, comp545minJ, comp2134minVal, comp2134minI, comp2134minJ);
    wire [11:0] comp2135minVal;
    wire [5:0] comp2135minI, comp2135minJ;
    Comparator comp2135(comp546minVal, comp546minI, comp546minJ, comp547minVal, comp547minI, comp547minJ, comp2135minVal, comp2135minI, comp2135minJ);
    wire [11:0] comp2136minVal;
    wire [5:0] comp2136minI, comp2136minJ;
    Comparator comp2136(comp548minVal, comp548minI, comp548minJ, comp549minVal, comp549minI, comp549minJ, comp2136minVal, comp2136minI, comp2136minJ);
    wire [11:0] comp2137minVal;
    wire [5:0] comp2137minI, comp2137minJ;
    Comparator comp2137(comp550minVal, comp550minI, comp550minJ, comp551minVal, comp551minI, comp551minJ, comp2137minVal, comp2137minI, comp2137minJ);
    wire [11:0] comp2138minVal;
    wire [5:0] comp2138minI, comp2138minJ;
    Comparator comp2138(comp552minVal, comp552minI, comp552minJ, comp553minVal, comp553minI, comp553minJ, comp2138minVal, comp2138minI, comp2138minJ);
    wire [11:0] comp2139minVal;
    wire [5:0] comp2139minI, comp2139minJ;
    Comparator comp2139(comp554minVal, comp554minI, comp554minJ, comp555minVal, comp555minI, comp555minJ, comp2139minVal, comp2139minI, comp2139minJ);
    wire [11:0] comp2140minVal;
    wire [5:0] comp2140minI, comp2140minJ;
    Comparator comp2140(comp556minVal, comp556minI, comp556minJ, comp557minVal, comp557minI, comp557minJ, comp2140minVal, comp2140minI, comp2140minJ);
    wire [11:0] comp2141minVal;
    wire [5:0] comp2141minI, comp2141minJ;
    Comparator comp2141(comp558minVal, comp558minI, comp558minJ, comp559minVal, comp559minI, comp559minJ, comp2141minVal, comp2141minI, comp2141minJ);
    wire [11:0] comp2142minVal;
    wire [5:0] comp2142minI, comp2142minJ;
    Comparator comp2142(comp560minVal, comp560minI, comp560minJ, comp561minVal, comp561minI, comp561minJ, comp2142minVal, comp2142minI, comp2142minJ);
    wire [11:0] comp2143minVal;
    wire [5:0] comp2143minI, comp2143minJ;
    Comparator comp2143(comp562minVal, comp562minI, comp562minJ, comp563minVal, comp563minI, comp563minJ, comp2143minVal, comp2143minI, comp2143minJ);
    wire [11:0] comp2144minVal;
    wire [5:0] comp2144minI, comp2144minJ;
    Comparator comp2144(comp564minVal, comp564minI, comp564minJ, comp565minVal, comp565minI, comp565minJ, comp2144minVal, comp2144minI, comp2144minJ);
    wire [11:0] comp2145minVal;
    wire [5:0] comp2145minI, comp2145minJ;
    Comparator comp2145(comp566minVal, comp566minI, comp566minJ, comp567minVal, comp567minI, comp567minJ, comp2145minVal, comp2145minI, comp2145minJ);
    wire [11:0] comp2146minVal;
    wire [5:0] comp2146minI, comp2146minJ;
    Comparator comp2146(comp568minVal, comp568minI, comp568minJ, comp569minVal, comp569minI, comp569minJ, comp2146minVal, comp2146minI, comp2146minJ);
    wire [11:0] comp2147minVal;
    wire [5:0] comp2147minI, comp2147minJ;
    Comparator comp2147(comp570minVal, comp570minI, comp570minJ, comp571minVal, comp571minI, comp571minJ, comp2147minVal, comp2147minI, comp2147minJ);
    wire [11:0] comp2148minVal;
    wire [5:0] comp2148minI, comp2148minJ;
    Comparator comp2148(comp572minVal, comp572minI, comp572minJ, comp573minVal, comp573minI, comp573minJ, comp2148minVal, comp2148minI, comp2148minJ);
    wire [11:0] comp2149minVal;
    wire [5:0] comp2149minI, comp2149minJ;
    Comparator comp2149(comp574minVal, comp574minI, comp574minJ, comp575minVal, comp575minI, comp575minJ, comp2149minVal, comp2149minI, comp2149minJ);
    wire [11:0] comp2150minVal;
    wire [5:0] comp2150minI, comp2150minJ;
    Comparator comp2150(comp576minVal, comp576minI, comp576minJ, comp577minVal, comp577minI, comp577minJ, comp2150minVal, comp2150minI, comp2150minJ);
    wire [11:0] comp2151minVal;
    wire [5:0] comp2151minI, comp2151minJ;
    Comparator comp2151(comp578minVal, comp578minI, comp578minJ, comp579minVal, comp579minI, comp579minJ, comp2151minVal, comp2151minI, comp2151minJ);
    wire [11:0] comp2152minVal;
    wire [5:0] comp2152minI, comp2152minJ;
    Comparator comp2152(comp580minVal, comp580minI, comp580minJ, comp581minVal, comp581minI, comp581minJ, comp2152minVal, comp2152minI, comp2152minJ);
    wire [11:0] comp2153minVal;
    wire [5:0] comp2153minI, comp2153minJ;
    Comparator comp2153(comp582minVal, comp582minI, comp582minJ, comp583minVal, comp583minI, comp583minJ, comp2153minVal, comp2153minI, comp2153minJ);
    wire [11:0] comp2154minVal;
    wire [5:0] comp2154minI, comp2154minJ;
    Comparator comp2154(comp584minVal, comp584minI, comp584minJ, comp585minVal, comp585minI, comp585minJ, comp2154minVal, comp2154minI, comp2154minJ);
    wire [11:0] comp2155minVal;
    wire [5:0] comp2155minI, comp2155minJ;
    Comparator comp2155(comp586minVal, comp586minI, comp586minJ, comp587minVal, comp587minI, comp587minJ, comp2155minVal, comp2155minI, comp2155minJ);
    wire [11:0] comp2156minVal;
    wire [5:0] comp2156minI, comp2156minJ;
    Comparator comp2156(comp588minVal, comp588minI, comp588minJ, comp589minVal, comp589minI, comp589minJ, comp2156minVal, comp2156minI, comp2156minJ);
    wire [11:0] comp2157minVal;
    wire [5:0] comp2157minI, comp2157minJ;
    Comparator comp2157(comp590minVal, comp590minI, comp590minJ, comp591minVal, comp591minI, comp591minJ, comp2157minVal, comp2157minI, comp2157minJ);
    wire [11:0] comp2158minVal;
    wire [5:0] comp2158minI, comp2158minJ;
    Comparator comp2158(comp592minVal, comp592minI, comp592minJ, comp593minVal, comp593minI, comp593minJ, comp2158minVal, comp2158minI, comp2158minJ);
    wire [11:0] comp2159minVal;
    wire [5:0] comp2159minI, comp2159minJ;
    Comparator comp2159(comp594minVal, comp594minI, comp594minJ, comp595minVal, comp595minI, comp595minJ, comp2159minVal, comp2159minI, comp2159minJ);
    wire [11:0] comp2160minVal;
    wire [5:0] comp2160minI, comp2160minJ;
    Comparator comp2160(comp596minVal, comp596minI, comp596minJ, comp597minVal, comp597minI, comp597minJ, comp2160minVal, comp2160minI, comp2160minJ);
    wire [11:0] comp2161minVal;
    wire [5:0] comp2161minI, comp2161minJ;
    Comparator comp2161(comp598minVal, comp598minI, comp598minJ, comp599minVal, comp599minI, comp599minJ, comp2161minVal, comp2161minI, comp2161minJ);
    wire [11:0] comp2162minVal;
    wire [5:0] comp2162minI, comp2162minJ;
    Comparator comp2162(comp600minVal, comp600minI, comp600minJ, comp601minVal, comp601minI, comp601minJ, comp2162minVal, comp2162minI, comp2162minJ);
    wire [11:0] comp2163minVal;
    wire [5:0] comp2163minI, comp2163minJ;
    Comparator comp2163(comp602minVal, comp602minI, comp602minJ, comp603minVal, comp603minI, comp603minJ, comp2163minVal, comp2163minI, comp2163minJ);
    wire [11:0] comp2164minVal;
    wire [5:0] comp2164minI, comp2164minJ;
    Comparator comp2164(comp604minVal, comp604minI, comp604minJ, comp605minVal, comp605minI, comp605minJ, comp2164minVal, comp2164minI, comp2164minJ);
    wire [11:0] comp2165minVal;
    wire [5:0] comp2165minI, comp2165minJ;
    Comparator comp2165(comp606minVal, comp606minI, comp606minJ, comp607minVal, comp607minI, comp607minJ, comp2165minVal, comp2165minI, comp2165minJ);
    wire [11:0] comp2166minVal;
    wire [5:0] comp2166minI, comp2166minJ;
    Comparator comp2166(comp608minVal, comp608minI, comp608minJ, comp609minVal, comp609minI, comp609minJ, comp2166minVal, comp2166minI, comp2166minJ);
    wire [11:0] comp2167minVal;
    wire [5:0] comp2167minI, comp2167minJ;
    Comparator comp2167(comp610minVal, comp610minI, comp610minJ, comp611minVal, comp611minI, comp611minJ, comp2167minVal, comp2167minI, comp2167minJ);
    wire [11:0] comp2168minVal;
    wire [5:0] comp2168minI, comp2168minJ;
    Comparator comp2168(comp612minVal, comp612minI, comp612minJ, comp613minVal, comp613minI, comp613minJ, comp2168minVal, comp2168minI, comp2168minJ);
    wire [11:0] comp2169minVal;
    wire [5:0] comp2169minI, comp2169minJ;
    Comparator comp2169(comp614minVal, comp614minI, comp614minJ, comp615minVal, comp615minI, comp615minJ, comp2169minVal, comp2169minI, comp2169minJ);
    wire [11:0] comp2170minVal;
    wire [5:0] comp2170minI, comp2170minJ;
    Comparator comp2170(comp616minVal, comp616minI, comp616minJ, comp617minVal, comp617minI, comp617minJ, comp2170minVal, comp2170minI, comp2170minJ);
    wire [11:0] comp2171minVal;
    wire [5:0] comp2171minI, comp2171minJ;
    Comparator comp2171(comp618minVal, comp618minI, comp618minJ, comp619minVal, comp619minI, comp619minJ, comp2171minVal, comp2171minI, comp2171minJ);
    wire [11:0] comp2172minVal;
    wire [5:0] comp2172minI, comp2172minJ;
    Comparator comp2172(comp620minVal, comp620minI, comp620minJ, comp621minVal, comp621minI, comp621minJ, comp2172minVal, comp2172minI, comp2172minJ);
    wire [11:0] comp2173minVal;
    wire [5:0] comp2173minI, comp2173minJ;
    Comparator comp2173(comp622minVal, comp622minI, comp622minJ, comp623minVal, comp623minI, comp623minJ, comp2173minVal, comp2173minI, comp2173minJ);
    wire [11:0] comp2174minVal;
    wire [5:0] comp2174minI, comp2174minJ;
    Comparator comp2174(comp624minVal, comp624minI, comp624minJ, comp625minVal, comp625minI, comp625minJ, comp2174minVal, comp2174minI, comp2174minJ);
    wire [11:0] comp2175minVal;
    wire [5:0] comp2175minI, comp2175minJ;
    Comparator comp2175(comp626minVal, comp626minI, comp626minJ, comp627minVal, comp627minI, comp627minJ, comp2175minVal, comp2175minI, comp2175minJ);
    wire [11:0] comp2176minVal;
    wire [5:0] comp2176minI, comp2176minJ;
    Comparator comp2176(comp628minVal, comp628minI, comp628minJ, comp629minVal, comp629minI, comp629minJ, comp2176minVal, comp2176minI, comp2176minJ);
    wire [11:0] comp2177minVal;
    wire [5:0] comp2177minI, comp2177minJ;
    Comparator comp2177(comp630minVal, comp630minI, comp630minJ, comp631minVal, comp631minI, comp631minJ, comp2177minVal, comp2177minI, comp2177minJ);
    wire [11:0] comp2178minVal;
    wire [5:0] comp2178minI, comp2178minJ;
    Comparator comp2178(comp632minVal, comp632minI, comp632minJ, comp633minVal, comp633minI, comp633minJ, comp2178minVal, comp2178minI, comp2178minJ);
    wire [11:0] comp2179minVal;
    wire [5:0] comp2179minI, comp2179minJ;
    Comparator comp2179(comp634minVal, comp634minI, comp634minJ, comp635minVal, comp635minI, comp635minJ, comp2179minVal, comp2179minI, comp2179minJ);
    wire [11:0] comp2180minVal;
    wire [5:0] comp2180minI, comp2180minJ;
    Comparator comp2180(comp636minVal, comp636minI, comp636minJ, comp637minVal, comp637minI, comp637minJ, comp2180minVal, comp2180minI, comp2180minJ);
    wire [11:0] comp2181minVal;
    wire [5:0] comp2181minI, comp2181minJ;
    Comparator comp2181(comp638minVal, comp638minI, comp638minJ, comp639minVal, comp639minI, comp639minJ, comp2181minVal, comp2181minI, comp2181minJ);
    wire [11:0] comp2182minVal;
    wire [5:0] comp2182minI, comp2182minJ;
    Comparator comp2182(comp640minVal, comp640minI, comp640minJ, comp641minVal, comp641minI, comp641minJ, comp2182minVal, comp2182minI, comp2182minJ);
    wire [11:0] comp2183minVal;
    wire [5:0] comp2183minI, comp2183minJ;
    Comparator comp2183(comp642minVal, comp642minI, comp642minJ, comp643minVal, comp643minI, comp643minJ, comp2183minVal, comp2183minI, comp2183minJ);
    wire [11:0] comp2184minVal;
    wire [5:0] comp2184minI, comp2184minJ;
    Comparator comp2184(comp644minVal, comp644minI, comp644minJ, comp645minVal, comp645minI, comp645minJ, comp2184minVal, comp2184minI, comp2184minJ);
    wire [11:0] comp2185minVal;
    wire [5:0] comp2185minI, comp2185minJ;
    Comparator comp2185(comp646minVal, comp646minI, comp646minJ, comp647minVal, comp647minI, comp647minJ, comp2185minVal, comp2185minI, comp2185minJ);
    wire [11:0] comp2186minVal;
    wire [5:0] comp2186minI, comp2186minJ;
    Comparator comp2186(comp648minVal, comp648minI, comp648minJ, comp649minVal, comp649minI, comp649minJ, comp2186minVal, comp2186minI, comp2186minJ);
    wire [11:0] comp2187minVal;
    wire [5:0] comp2187minI, comp2187minJ;
    Comparator comp2187(comp650minVal, comp650minI, comp650minJ, comp651minVal, comp651minI, comp651minJ, comp2187minVal, comp2187minI, comp2187minJ);
    wire [11:0] comp2188minVal;
    wire [5:0] comp2188minI, comp2188minJ;
    Comparator comp2188(comp652minVal, comp652minI, comp652minJ, comp653minVal, comp653minI, comp653minJ, comp2188minVal, comp2188minI, comp2188minJ);
    wire [11:0] comp2189minVal;
    wire [5:0] comp2189minI, comp2189minJ;
    Comparator comp2189(comp654minVal, comp654minI, comp654minJ, comp655minVal, comp655minI, comp655minJ, comp2189minVal, comp2189minI, comp2189minJ);
    wire [11:0] comp2190minVal;
    wire [5:0] comp2190minI, comp2190minJ;
    Comparator comp2190(comp656minVal, comp656minI, comp656minJ, comp657minVal, comp657minI, comp657minJ, comp2190minVal, comp2190minI, comp2190minJ);
    wire [11:0] comp2191minVal;
    wire [5:0] comp2191minI, comp2191minJ;
    Comparator comp2191(comp658minVal, comp658minI, comp658minJ, comp659minVal, comp659minI, comp659minJ, comp2191minVal, comp2191minI, comp2191minJ);
    wire [11:0] comp2192minVal;
    wire [5:0] comp2192minI, comp2192minJ;
    Comparator comp2192(comp660minVal, comp660minI, comp660minJ, comp661minVal, comp661minI, comp661minJ, comp2192minVal, comp2192minI, comp2192minJ);
    wire [11:0] comp2193minVal;
    wire [5:0] comp2193minI, comp2193minJ;
    Comparator comp2193(comp662minVal, comp662minI, comp662minJ, comp663minVal, comp663minI, comp663minJ, comp2193minVal, comp2193minI, comp2193minJ);
    wire [11:0] comp2194minVal;
    wire [5:0] comp2194minI, comp2194minJ;
    Comparator comp2194(comp664minVal, comp664minI, comp664minJ, comp665minVal, comp665minI, comp665minJ, comp2194minVal, comp2194minI, comp2194minJ);
    wire [11:0] comp2195minVal;
    wire [5:0] comp2195minI, comp2195minJ;
    Comparator comp2195(comp666minVal, comp666minI, comp666minJ, comp667minVal, comp667minI, comp667minJ, comp2195minVal, comp2195minI, comp2195minJ);
    wire [11:0] comp2196minVal;
    wire [5:0] comp2196minI, comp2196minJ;
    Comparator comp2196(comp668minVal, comp668minI, comp668minJ, comp669minVal, comp669minI, comp669minJ, comp2196minVal, comp2196minI, comp2196minJ);
    wire [11:0] comp2197minVal;
    wire [5:0] comp2197minI, comp2197minJ;
    Comparator comp2197(comp670minVal, comp670minI, comp670minJ, comp671minVal, comp671minI, comp671minJ, comp2197minVal, comp2197minI, comp2197minJ);
    wire [11:0] comp2198minVal;
    wire [5:0] comp2198minI, comp2198minJ;
    Comparator comp2198(comp672minVal, comp672minI, comp672minJ, comp673minVal, comp673minI, comp673minJ, comp2198minVal, comp2198minI, comp2198minJ);
    wire [11:0] comp2199minVal;
    wire [5:0] comp2199minI, comp2199minJ;
    Comparator comp2199(comp674minVal, comp674minI, comp674minJ, comp675minVal, comp675minI, comp675minJ, comp2199minVal, comp2199minI, comp2199minJ);
    wire [11:0] comp2200minVal;
    wire [5:0] comp2200minI, comp2200minJ;
    Comparator comp2200(comp676minVal, comp676minI, comp676minJ, comp677minVal, comp677minI, comp677minJ, comp2200minVal, comp2200minI, comp2200minJ);
    wire [11:0] comp2201minVal;
    wire [5:0] comp2201minI, comp2201minJ;
    Comparator comp2201(comp678minVal, comp678minI, comp678minJ, comp679minVal, comp679minI, comp679minJ, comp2201minVal, comp2201minI, comp2201minJ);
    wire [11:0] comp2202minVal;
    wire [5:0] comp2202minI, comp2202minJ;
    Comparator comp2202(comp680minVal, comp680minI, comp680minJ, comp681minVal, comp681minI, comp681minJ, comp2202minVal, comp2202minI, comp2202minJ);
    wire [11:0] comp2203minVal;
    wire [5:0] comp2203minI, comp2203minJ;
    Comparator comp2203(comp682minVal, comp682minI, comp682minJ, comp683minVal, comp683minI, comp683minJ, comp2203minVal, comp2203minI, comp2203minJ);
    wire [11:0] comp2204minVal;
    wire [5:0] comp2204minI, comp2204minJ;
    Comparator comp2204(comp684minVal, comp684minI, comp684minJ, comp685minVal, comp685minI, comp685minJ, comp2204minVal, comp2204minI, comp2204minJ);
    wire [11:0] comp2205minVal;
    wire [5:0] comp2205minI, comp2205minJ;
    Comparator comp2205(comp686minVal, comp686minI, comp686minJ, comp687minVal, comp687minI, comp687minJ, comp2205minVal, comp2205minI, comp2205minJ);
    wire [11:0] comp2206minVal;
    wire [5:0] comp2206minI, comp2206minJ;
    Comparator comp2206(comp688minVal, comp688minI, comp688minJ, comp689minVal, comp689minI, comp689minJ, comp2206minVal, comp2206minI, comp2206minJ);
    wire [11:0] comp2207minVal;
    wire [5:0] comp2207minI, comp2207minJ;
    Comparator comp2207(comp690minVal, comp690minI, comp690minJ, comp691minVal, comp691minI, comp691minJ, comp2207minVal, comp2207minI, comp2207minJ);
    wire [11:0] comp2208minVal;
    wire [5:0] comp2208minI, comp2208minJ;
    Comparator comp2208(comp692minVal, comp692minI, comp692minJ, comp693minVal, comp693minI, comp693minJ, comp2208minVal, comp2208minI, comp2208minJ);
    wire [11:0] comp2209minVal;
    wire [5:0] comp2209minI, comp2209minJ;
    Comparator comp2209(comp694minVal, comp694minI, comp694minJ, comp695minVal, comp695minI, comp695minJ, comp2209minVal, comp2209minI, comp2209minJ);
    wire [11:0] comp2210minVal;
    wire [5:0] comp2210minI, comp2210minJ;
    Comparator comp2210(comp696minVal, comp696minI, comp696minJ, comp697minVal, comp697minI, comp697minJ, comp2210minVal, comp2210minI, comp2210minJ);
    wire [11:0] comp2211minVal;
    wire [5:0] comp2211minI, comp2211minJ;
    Comparator comp2211(comp698minVal, comp698minI, comp698minJ, comp699minVal, comp699minI, comp699minJ, comp2211minVal, comp2211minI, comp2211minJ);
    wire [11:0] comp2212minVal;
    wire [5:0] comp2212minI, comp2212minJ;
    Comparator comp2212(comp700minVal, comp700minI, comp700minJ, comp701minVal, comp701minI, comp701minJ, comp2212minVal, comp2212minI, comp2212minJ);
    wire [11:0] comp2213minVal;
    wire [5:0] comp2213minI, comp2213minJ;
    Comparator comp2213(comp702minVal, comp702minI, comp702minJ, comp703minVal, comp703minI, comp703minJ, comp2213minVal, comp2213minI, comp2213minJ);
    wire [11:0] comp2214minVal;
    wire [5:0] comp2214minI, comp2214minJ;
    Comparator comp2214(comp704minVal, comp704minI, comp704minJ, comp705minVal, comp705minI, comp705minJ, comp2214minVal, comp2214minI, comp2214minJ);
    wire [11:0] comp2215minVal;
    wire [5:0] comp2215minI, comp2215minJ;
    Comparator comp2215(comp706minVal, comp706minI, comp706minJ, comp707minVal, comp707minI, comp707minJ, comp2215minVal, comp2215minI, comp2215minJ);
    wire [11:0] comp2216minVal;
    wire [5:0] comp2216minI, comp2216minJ;
    Comparator comp2216(comp708minVal, comp708minI, comp708minJ, comp709minVal, comp709minI, comp709minJ, comp2216minVal, comp2216minI, comp2216minJ);
    wire [11:0] comp2217minVal;
    wire [5:0] comp2217minI, comp2217minJ;
    Comparator comp2217(comp710minVal, comp710minI, comp710minJ, comp711minVal, comp711minI, comp711minJ, comp2217minVal, comp2217minI, comp2217minJ);
    wire [11:0] comp2218minVal;
    wire [5:0] comp2218minI, comp2218minJ;
    Comparator comp2218(comp712minVal, comp712minI, comp712minJ, comp713minVal, comp713minI, comp713minJ, comp2218minVal, comp2218minI, comp2218minJ);
    wire [11:0] comp2219minVal;
    wire [5:0] comp2219minI, comp2219minJ;
    Comparator comp2219(comp714minVal, comp714minI, comp714minJ, comp715minVal, comp715minI, comp715minJ, comp2219minVal, comp2219minI, comp2219minJ);
    wire [11:0] comp2220minVal;
    wire [5:0] comp2220minI, comp2220minJ;
    Comparator comp2220(comp716minVal, comp716minI, comp716minJ, comp717minVal, comp717minI, comp717minJ, comp2220minVal, comp2220minI, comp2220minJ);
    wire [11:0] comp2221minVal;
    wire [5:0] comp2221minI, comp2221minJ;
    Comparator comp2221(comp718minVal, comp718minI, comp718minJ, comp719minVal, comp719minI, comp719minJ, comp2221minVal, comp2221minI, comp2221minJ);
    wire [11:0] comp2222minVal;
    wire [5:0] comp2222minI, comp2222minJ;
    Comparator comp2222(comp720minVal, comp720minI, comp720minJ, comp721minVal, comp721minI, comp721minJ, comp2222minVal, comp2222minI, comp2222minJ);
    wire [11:0] comp2223minVal;
    wire [5:0] comp2223minI, comp2223minJ;
    Comparator comp2223(comp722minVal, comp722minI, comp722minJ, comp723minVal, comp723minI, comp723minJ, comp2223minVal, comp2223minI, comp2223minJ);
    wire [11:0] comp2224minVal;
    wire [5:0] comp2224minI, comp2224minJ;
    Comparator comp2224(comp724minVal, comp724minI, comp724minJ, comp725minVal, comp725minI, comp725minJ, comp2224minVal, comp2224minI, comp2224minJ);
    wire [11:0] comp2225minVal;
    wire [5:0] comp2225minI, comp2225minJ;
    Comparator comp2225(comp726minVal, comp726minI, comp726minJ, comp727minVal, comp727minI, comp727minJ, comp2225minVal, comp2225minI, comp2225minJ);
    wire [11:0] comp2226minVal;
    wire [5:0] comp2226minI, comp2226minJ;
    Comparator comp2226(comp728minVal, comp728minI, comp728minJ, comp729minVal, comp729minI, comp729minJ, comp2226minVal, comp2226minI, comp2226minJ);
    wire [11:0] comp2227minVal;
    wire [5:0] comp2227minI, comp2227minJ;
    Comparator comp2227(comp730minVal, comp730minI, comp730minJ, comp731minVal, comp731minI, comp731minJ, comp2227minVal, comp2227minI, comp2227minJ);
    wire [11:0] comp2228minVal;
    wire [5:0] comp2228minI, comp2228minJ;
    Comparator comp2228(comp732minVal, comp732minI, comp732minJ, comp733minVal, comp733minI, comp733minJ, comp2228minVal, comp2228minI, comp2228minJ);
    wire [11:0] comp2229minVal;
    wire [5:0] comp2229minI, comp2229minJ;
    Comparator comp2229(comp734minVal, comp734minI, comp734minJ, comp735minVal, comp735minI, comp735minJ, comp2229minVal, comp2229minI, comp2229minJ);
    wire [11:0] comp2230minVal;
    wire [5:0] comp2230minI, comp2230minJ;
    Comparator comp2230(comp736minVal, comp736minI, comp736minJ, comp737minVal, comp737minI, comp737minJ, comp2230minVal, comp2230minI, comp2230minJ);
    wire [11:0] comp2231minVal;
    wire [5:0] comp2231minI, comp2231minJ;
    Comparator comp2231(comp738minVal, comp738minI, comp738minJ, comp739minVal, comp739minI, comp739minJ, comp2231minVal, comp2231minI, comp2231minJ);
    wire [11:0] comp2232minVal;
    wire [5:0] comp2232minI, comp2232minJ;
    Comparator comp2232(comp740minVal, comp740minI, comp740minJ, comp741minVal, comp741minI, comp741minJ, comp2232minVal, comp2232minI, comp2232minJ);
    wire [11:0] comp2233minVal;
    wire [5:0] comp2233minI, comp2233minJ;
    Comparator comp2233(comp742minVal, comp742minI, comp742minJ, comp743minVal, comp743minI, comp743minJ, comp2233minVal, comp2233minI, comp2233minJ);
    wire [11:0] comp2234minVal;
    wire [5:0] comp2234minI, comp2234minJ;
    Comparator comp2234(comp744minVal, comp744minI, comp744minJ, comp745minVal, comp745minI, comp745minJ, comp2234minVal, comp2234minI, comp2234minJ);
    wire [11:0] comp2235minVal;
    wire [5:0] comp2235minI, comp2235minJ;
    Comparator comp2235(comp746minVal, comp746minI, comp746minJ, comp747minVal, comp747minI, comp747minJ, comp2235minVal, comp2235minI, comp2235minJ);
    wire [11:0] comp2236minVal;
    wire [5:0] comp2236minI, comp2236minJ;
    Comparator comp2236(comp748minVal, comp748minI, comp748minJ, comp749minVal, comp749minI, comp749minJ, comp2236minVal, comp2236minI, comp2236minJ);
    wire [11:0] comp2237minVal;
    wire [5:0] comp2237minI, comp2237minJ;
    Comparator comp2237(comp750minVal, comp750minI, comp750minJ, comp751minVal, comp751minI, comp751minJ, comp2237minVal, comp2237minI, comp2237minJ);
    wire [11:0] comp2238minVal;
    wire [5:0] comp2238minI, comp2238minJ;
    Comparator comp2238(comp752minVal, comp752minI, comp752minJ, comp753minVal, comp753minI, comp753minJ, comp2238minVal, comp2238minI, comp2238minJ);
    wire [11:0] comp2239minVal;
    wire [5:0] comp2239minI, comp2239minJ;
    Comparator comp2239(comp754minVal, comp754minI, comp754minJ, comp755minVal, comp755minI, comp755minJ, comp2239minVal, comp2239minI, comp2239minJ);
    wire [11:0] comp2240minVal;
    wire [5:0] comp2240minI, comp2240minJ;
    Comparator comp2240(comp756minVal, comp756minI, comp756minJ, comp757minVal, comp757minI, comp757minJ, comp2240minVal, comp2240minI, comp2240minJ);
    wire [11:0] comp2241minVal;
    wire [5:0] comp2241minI, comp2241minJ;
    Comparator comp2241(comp758minVal, comp758minI, comp758minJ, comp759minVal, comp759minI, comp759minJ, comp2241minVal, comp2241minI, comp2241minJ);
    wire [11:0] comp2242minVal;
    wire [5:0] comp2242minI, comp2242minJ;
    Comparator comp2242(comp760minVal, comp760minI, comp760minJ, comp761minVal, comp761minI, comp761minJ, comp2242minVal, comp2242minI, comp2242minJ);
    wire [11:0] comp2243minVal;
    wire [5:0] comp2243minI, comp2243minJ;
    Comparator comp2243(comp762minVal, comp762minI, comp762minJ, comp763minVal, comp763minI, comp763minJ, comp2243minVal, comp2243minI, comp2243minJ);
    wire [11:0] comp2244minVal;
    wire [5:0] comp2244minI, comp2244minJ;
    Comparator comp2244(comp764minVal, comp764minI, comp764minJ, comp765minVal, comp765minI, comp765minJ, comp2244minVal, comp2244minI, comp2244minJ);
    wire [11:0] comp2245minVal;
    wire [5:0] comp2245minI, comp2245minJ;
    Comparator comp2245(comp766minVal, comp766minI, comp766minJ, comp767minVal, comp767minI, comp767minJ, comp2245minVal, comp2245minI, comp2245minJ);
    wire [11:0] comp2246minVal;
    wire [5:0] comp2246minI, comp2246minJ;
    Comparator comp2246(comp768minVal, comp768minI, comp768minJ, comp769minVal, comp769minI, comp769minJ, comp2246minVal, comp2246minI, comp2246minJ);
    wire [11:0] comp2247minVal;
    wire [5:0] comp2247minI, comp2247minJ;
    Comparator comp2247(comp770minVal, comp770minI, comp770minJ, comp771minVal, comp771minI, comp771minJ, comp2247minVal, comp2247minI, comp2247minJ);
    wire [11:0] comp2248minVal;
    wire [5:0] comp2248minI, comp2248minJ;
    Comparator comp2248(comp772minVal, comp772minI, comp772minJ, comp773minVal, comp773minI, comp773minJ, comp2248minVal, comp2248minI, comp2248minJ);
    wire [11:0] comp2249minVal;
    wire [5:0] comp2249minI, comp2249minJ;
    Comparator comp2249(comp774minVal, comp774minI, comp774minJ, comp775minVal, comp775minI, comp775minJ, comp2249minVal, comp2249minI, comp2249minJ);
    wire [11:0] comp2250minVal;
    wire [5:0] comp2250minI, comp2250minJ;
    Comparator comp2250(comp776minVal, comp776minI, comp776minJ, comp777minVal, comp777minI, comp777minJ, comp2250minVal, comp2250minI, comp2250minJ);
    wire [11:0] comp2251minVal;
    wire [5:0] comp2251minI, comp2251minJ;
    Comparator comp2251(comp778minVal, comp778minI, comp778minJ, comp779minVal, comp779minI, comp779minJ, comp2251minVal, comp2251minI, comp2251minJ);
    wire [11:0] comp2252minVal;
    wire [5:0] comp2252minI, comp2252minJ;
    Comparator comp2252(comp780minVal, comp780minI, comp780minJ, comp781minVal, comp781minI, comp781minJ, comp2252minVal, comp2252minI, comp2252minJ);
    wire [11:0] comp2253minVal;
    wire [5:0] comp2253minI, comp2253minJ;
    Comparator comp2253(comp782minVal, comp782minI, comp782minJ, comp783minVal, comp783minI, comp783minJ, comp2253minVal, comp2253minI, comp2253minJ);
    wire [11:0] comp2254minVal;
    wire [5:0] comp2254minI, comp2254minJ;
    Comparator comp2254(comp784minVal, comp784minI, comp784minJ, comp785minVal, comp785minI, comp785minJ, comp2254minVal, comp2254minI, comp2254minJ);
    wire [11:0] comp2255minVal;
    wire [5:0] comp2255minI, comp2255minJ;
    Comparator comp2255(comp786minVal, comp786minI, comp786minJ, comp787minVal, comp787minI, comp787minJ, comp2255minVal, comp2255minI, comp2255minJ);
    wire [11:0] comp2256minVal;
    wire [5:0] comp2256minI, comp2256minJ;
    Comparator comp2256(comp788minVal, comp788minI, comp788minJ, comp789minVal, comp789minI, comp789minJ, comp2256minVal, comp2256minI, comp2256minJ);
    wire [11:0] comp2257minVal;
    wire [5:0] comp2257minI, comp2257minJ;
    Comparator comp2257(comp790minVal, comp790minI, comp790minJ, comp791minVal, comp791minI, comp791minJ, comp2257minVal, comp2257minI, comp2257minJ);
    wire [11:0] comp2258minVal;
    wire [5:0] comp2258minI, comp2258minJ;
    Comparator comp2258(comp792minVal, comp792minI, comp792minJ, comp793minVal, comp793minI, comp793minJ, comp2258minVal, comp2258minI, comp2258minJ);
    wire [11:0] comp2259minVal;
    wire [5:0] comp2259minI, comp2259minJ;
    Comparator comp2259(comp794minVal, comp794minI, comp794minJ, comp795minVal, comp795minI, comp795minJ, comp2259minVal, comp2259minI, comp2259minJ);
    wire [11:0] comp2260minVal;
    wire [5:0] comp2260minI, comp2260minJ;
    Comparator comp2260(comp796minVal, comp796minI, comp796minJ, comp797minVal, comp797minI, comp797minJ, comp2260minVal, comp2260minI, comp2260minJ);
    wire [11:0] comp2261minVal;
    wire [5:0] comp2261minI, comp2261minJ;
    Comparator comp2261(comp798minVal, comp798minI, comp798minJ, comp799minVal, comp799minI, comp799minJ, comp2261minVal, comp2261minI, comp2261minJ);
    wire [11:0] comp2262minVal;
    wire [5:0] comp2262minI, comp2262minJ;
    Comparator comp2262(comp800minVal, comp800minI, comp800minJ, comp801minVal, comp801minI, comp801minJ, comp2262minVal, comp2262minI, comp2262minJ);
    wire [11:0] comp2263minVal;
    wire [5:0] comp2263minI, comp2263minJ;
    Comparator comp2263(comp802minVal, comp802minI, comp802minJ, comp803minVal, comp803minI, comp803minJ, comp2263minVal, comp2263minI, comp2263minJ);
    wire [11:0] comp2264minVal;
    wire [5:0] comp2264minI, comp2264minJ;
    Comparator comp2264(comp804minVal, comp804minI, comp804minJ, comp805minVal, comp805minI, comp805minJ, comp2264minVal, comp2264minI, comp2264minJ);
    wire [11:0] comp2265minVal;
    wire [5:0] comp2265minI, comp2265minJ;
    Comparator comp2265(comp806minVal, comp806minI, comp806minJ, comp807minVal, comp807minI, comp807minJ, comp2265minVal, comp2265minI, comp2265minJ);
    wire [11:0] comp2266minVal;
    wire [5:0] comp2266minI, comp2266minJ;
    Comparator comp2266(comp808minVal, comp808minI, comp808minJ, comp809minVal, comp809minI, comp809minJ, comp2266minVal, comp2266minI, comp2266minJ);
    wire [11:0] comp2267minVal;
    wire [5:0] comp2267minI, comp2267minJ;
    Comparator comp2267(comp810minVal, comp810minI, comp810minJ, comp811minVal, comp811minI, comp811minJ, comp2267minVal, comp2267minI, comp2267minJ);
    wire [11:0] comp2268minVal;
    wire [5:0] comp2268minI, comp2268minJ;
    Comparator comp2268(comp812minVal, comp812minI, comp812minJ, comp813minVal, comp813minI, comp813minJ, comp2268minVal, comp2268minI, comp2268minJ);
    wire [11:0] comp2269minVal;
    wire [5:0] comp2269minI, comp2269minJ;
    Comparator comp2269(comp814minVal, comp814minI, comp814minJ, comp815minVal, comp815minI, comp815minJ, comp2269minVal, comp2269minI, comp2269minJ);
    wire [11:0] comp2270minVal;
    wire [5:0] comp2270minI, comp2270minJ;
    Comparator comp2270(comp816minVal, comp816minI, comp816minJ, comp817minVal, comp817minI, comp817minJ, comp2270minVal, comp2270minI, comp2270minJ);
    wire [11:0] comp2271minVal;
    wire [5:0] comp2271minI, comp2271minJ;
    Comparator comp2271(comp818minVal, comp818minI, comp818minJ, comp819minVal, comp819minI, comp819minJ, comp2271minVal, comp2271minI, comp2271minJ);
    wire [11:0] comp2272minVal;
    wire [5:0] comp2272minI, comp2272minJ;
    Comparator comp2272(comp820minVal, comp820minI, comp820minJ, comp821minVal, comp821minI, comp821minJ, comp2272minVal, comp2272minI, comp2272minJ);
    wire [11:0] comp2273minVal;
    wire [5:0] comp2273minI, comp2273minJ;
    Comparator comp2273(comp822minVal, comp822minI, comp822minJ, comp823minVal, comp823minI, comp823minJ, comp2273minVal, comp2273minI, comp2273minJ);
    wire [11:0] comp2274minVal;
    wire [5:0] comp2274minI, comp2274minJ;
    Comparator comp2274(comp824minVal, comp824minI, comp824minJ, comp825minVal, comp825minI, comp825minJ, comp2274minVal, comp2274minI, comp2274minJ);
    wire [11:0] comp2275minVal;
    wire [5:0] comp2275minI, comp2275minJ;
    Comparator comp2275(comp826minVal, comp826minI, comp826minJ, comp827minVal, comp827minI, comp827minJ, comp2275minVal, comp2275minI, comp2275minJ);
    wire [11:0] comp2276minVal;
    wire [5:0] comp2276minI, comp2276minJ;
    Comparator comp2276(comp828minVal, comp828minI, comp828minJ, comp829minVal, comp829minI, comp829minJ, comp2276minVal, comp2276minI, comp2276minJ);
    wire [11:0] comp2277minVal;
    wire [5:0] comp2277minI, comp2277minJ;
    Comparator comp2277(comp830minVal, comp830minI, comp830minJ, comp831minVal, comp831minI, comp831minJ, comp2277minVal, comp2277minI, comp2277minJ);
    wire [11:0] comp2278minVal;
    wire [5:0] comp2278minI, comp2278minJ;
    Comparator comp2278(comp832minVal, comp832minI, comp832minJ, comp833minVal, comp833minI, comp833minJ, comp2278minVal, comp2278minI, comp2278minJ);
    wire [11:0] comp2279minVal;
    wire [5:0] comp2279minI, comp2279minJ;
    Comparator comp2279(comp834minVal, comp834minI, comp834minJ, comp835minVal, comp835minI, comp835minJ, comp2279minVal, comp2279minI, comp2279minJ);
    wire [11:0] comp2280minVal;
    wire [5:0] comp2280minI, comp2280minJ;
    Comparator comp2280(comp836minVal, comp836minI, comp836minJ, comp837minVal, comp837minI, comp837minJ, comp2280minVal, comp2280minI, comp2280minJ);
    wire [11:0] comp2281minVal;
    wire [5:0] comp2281minI, comp2281minJ;
    Comparator comp2281(comp838minVal, comp838minI, comp838minJ, comp839minVal, comp839minI, comp839minJ, comp2281minVal, comp2281minI, comp2281minJ);
    wire [11:0] comp2282minVal;
    wire [5:0] comp2282minI, comp2282minJ;
    Comparator comp2282(comp840minVal, comp840minI, comp840minJ, comp841minVal, comp841minI, comp841minJ, comp2282minVal, comp2282minI, comp2282minJ);
    wire [11:0] comp2283minVal;
    wire [5:0] comp2283minI, comp2283minJ;
    Comparator comp2283(comp842minVal, comp842minI, comp842minJ, comp843minVal, comp843minI, comp843minJ, comp2283minVal, comp2283minI, comp2283minJ);
    wire [11:0] comp2284minVal;
    wire [5:0] comp2284minI, comp2284minJ;
    Comparator comp2284(comp844minVal, comp844minI, comp844minJ, comp845minVal, comp845minI, comp845minJ, comp2284minVal, comp2284minI, comp2284minJ);
    wire [11:0] comp2285minVal;
    wire [5:0] comp2285minI, comp2285minJ;
    Comparator comp2285(comp846minVal, comp846minI, comp846minJ, comp847minVal, comp847minI, comp847minJ, comp2285minVal, comp2285minI, comp2285minJ);
    wire [11:0] comp2286minVal;
    wire [5:0] comp2286minI, comp2286minJ;
    Comparator comp2286(comp848minVal, comp848minI, comp848minJ, comp849minVal, comp849minI, comp849minJ, comp2286minVal, comp2286minI, comp2286minJ);
    wire [11:0] comp2287minVal;
    wire [5:0] comp2287minI, comp2287minJ;
    Comparator comp2287(comp850minVal, comp850minI, comp850minJ, comp851minVal, comp851minI, comp851minJ, comp2287minVal, comp2287minI, comp2287minJ);
    wire [11:0] comp2288minVal;
    wire [5:0] comp2288minI, comp2288minJ;
    Comparator comp2288(comp852minVal, comp852minI, comp852minJ, comp853minVal, comp853minI, comp853minJ, comp2288minVal, comp2288minI, comp2288minJ);
    wire [11:0] comp2289minVal;
    wire [5:0] comp2289minI, comp2289minJ;
    Comparator comp2289(comp854minVal, comp854minI, comp854minJ, comp855minVal, comp855minI, comp855minJ, comp2289minVal, comp2289minI, comp2289minJ);
    wire [11:0] comp2290minVal;
    wire [5:0] comp2290minI, comp2290minJ;
    Comparator comp2290(comp856minVal, comp856minI, comp856minJ, comp857minVal, comp857minI, comp857minJ, comp2290minVal, comp2290minI, comp2290minJ);
    wire [11:0] comp2291minVal;
    wire [5:0] comp2291minI, comp2291minJ;
    Comparator comp2291(comp858minVal, comp858minI, comp858minJ, comp859minVal, comp859minI, comp859minJ, comp2291minVal, comp2291minI, comp2291minJ);
    wire [11:0] comp2292minVal;
    wire [5:0] comp2292minI, comp2292minJ;
    Comparator comp2292(comp860minVal, comp860minI, comp860minJ, comp861minVal, comp861minI, comp861minJ, comp2292minVal, comp2292minI, comp2292minJ);
    wire [11:0] comp2293minVal;
    wire [5:0] comp2293minI, comp2293minJ;
    Comparator comp2293(comp862minVal, comp862minI, comp862minJ, comp863minVal, comp863minI, comp863minJ, comp2293minVal, comp2293minI, comp2293minJ);
    wire [11:0] comp2294minVal;
    wire [5:0] comp2294minI, comp2294minJ;
    Comparator comp2294(comp864minVal, comp864minI, comp864minJ, comp865minVal, comp865minI, comp865minJ, comp2294minVal, comp2294minI, comp2294minJ);
    wire [11:0] comp2295minVal;
    wire [5:0] comp2295minI, comp2295minJ;
    Comparator comp2295(comp866minVal, comp866minI, comp866minJ, comp867minVal, comp867minI, comp867minJ, comp2295minVal, comp2295minI, comp2295minJ);
    wire [11:0] comp2296minVal;
    wire [5:0] comp2296minI, comp2296minJ;
    Comparator comp2296(comp868minVal, comp868minI, comp868minJ, comp869minVal, comp869minI, comp869minJ, comp2296minVal, comp2296minI, comp2296minJ);
    wire [11:0] comp2297minVal;
    wire [5:0] comp2297minI, comp2297minJ;
    Comparator comp2297(comp870minVal, comp870minI, comp870minJ, comp871minVal, comp871minI, comp871minJ, comp2297minVal, comp2297minI, comp2297minJ);
    wire [11:0] comp2298minVal;
    wire [5:0] comp2298minI, comp2298minJ;
    Comparator comp2298(comp872minVal, comp872minI, comp872minJ, comp873minVal, comp873minI, comp873minJ, comp2298minVal, comp2298minI, comp2298minJ);
    wire [11:0] comp2299minVal;
    wire [5:0] comp2299minI, comp2299minJ;
    Comparator comp2299(comp874minVal, comp874minI, comp874minJ, comp875minVal, comp875minI, comp875minJ, comp2299minVal, comp2299minI, comp2299minJ);
    wire [11:0] comp2300minVal;
    wire [5:0] comp2300minI, comp2300minJ;
    Comparator comp2300(comp876minVal, comp876minI, comp876minJ, comp877minVal, comp877minI, comp877minJ, comp2300minVal, comp2300minI, comp2300minJ);
    wire [11:0] comp2301minVal;
    wire [5:0] comp2301minI, comp2301minJ;
    Comparator comp2301(comp878minVal, comp878minI, comp878minJ, comp879minVal, comp879minI, comp879minJ, comp2301minVal, comp2301minI, comp2301minJ);
    wire [11:0] comp2302minVal;
    wire [5:0] comp2302minI, comp2302minJ;
    Comparator comp2302(comp880minVal, comp880minI, comp880minJ, comp881minVal, comp881minI, comp881minJ, comp2302minVal, comp2302minI, comp2302minJ);
    wire [11:0] comp2303minVal;
    wire [5:0] comp2303minI, comp2303minJ;
    Comparator comp2303(comp882minVal, comp882minI, comp882minJ, comp883minVal, comp883minI, comp883minJ, comp2303minVal, comp2303minI, comp2303minJ);
    wire [11:0] comp2304minVal;
    wire [5:0] comp2304minI, comp2304minJ;
    Comparator comp2304(comp884minVal, comp884minI, comp884minJ, comp885minVal, comp885minI, comp885minJ, comp2304minVal, comp2304minI, comp2304minJ);
    wire [11:0] comp2305minVal;
    wire [5:0] comp2305minI, comp2305minJ;
    Comparator comp2305(comp886minVal, comp886minI, comp886minJ, comp887minVal, comp887minI, comp887minJ, comp2305minVal, comp2305minI, comp2305minJ);
    wire [11:0] comp2306minVal;
    wire [5:0] comp2306minI, comp2306minJ;
    Comparator comp2306(comp888minVal, comp888minI, comp888minJ, comp889minVal, comp889minI, comp889minJ, comp2306minVal, comp2306minI, comp2306minJ);
    wire [11:0] comp2307minVal;
    wire [5:0] comp2307minI, comp2307minJ;
    Comparator comp2307(comp890minVal, comp890minI, comp890minJ, comp891minVal, comp891minI, comp891minJ, comp2307minVal, comp2307minI, comp2307minJ);
    wire [11:0] comp2308minVal;
    wire [5:0] comp2308minI, comp2308minJ;
    Comparator comp2308(comp892minVal, comp892minI, comp892minJ, comp893minVal, comp893minI, comp893minJ, comp2308minVal, comp2308minI, comp2308minJ);
    wire [11:0] comp2309minVal;
    wire [5:0] comp2309minI, comp2309minJ;
    Comparator comp2309(comp894minVal, comp894minI, comp894minJ, comp895minVal, comp895minI, comp895minJ, comp2309minVal, comp2309minI, comp2309minJ);
    wire [11:0] comp2310minVal;
    wire [5:0] comp2310minI, comp2310minJ;
    Comparator comp2310(comp896minVal, comp896minI, comp896minJ, comp897minVal, comp897minI, comp897minJ, comp2310minVal, comp2310minI, comp2310minJ);
    wire [11:0] comp2311minVal;
    wire [5:0] comp2311minI, comp2311minJ;
    Comparator comp2311(comp898minVal, comp898minI, comp898minJ, comp899minVal, comp899minI, comp899minJ, comp2311minVal, comp2311minI, comp2311minJ);
    wire [11:0] comp2312minVal;
    wire [5:0] comp2312minI, comp2312minJ;
    Comparator comp2312(comp900minVal, comp900minI, comp900minJ, comp901minVal, comp901minI, comp901minJ, comp2312minVal, comp2312minI, comp2312minJ);
    wire [11:0] comp2313minVal;
    wire [5:0] comp2313minI, comp2313minJ;
    Comparator comp2313(comp902minVal, comp902minI, comp902minJ, comp903minVal, comp903minI, comp903minJ, comp2313minVal, comp2313minI, comp2313minJ);
    wire [11:0] comp2314minVal;
    wire [5:0] comp2314minI, comp2314minJ;
    Comparator comp2314(comp904minVal, comp904minI, comp904minJ, comp905minVal, comp905minI, comp905minJ, comp2314minVal, comp2314minI, comp2314minJ);
    wire [11:0] comp2315minVal;
    wire [5:0] comp2315minI, comp2315minJ;
    Comparator comp2315(comp906minVal, comp906minI, comp906minJ, comp907minVal, comp907minI, comp907minJ, comp2315minVal, comp2315minI, comp2315minJ);
    wire [11:0] comp2316minVal;
    wire [5:0] comp2316minI, comp2316minJ;
    Comparator comp2316(comp908minVal, comp908minI, comp908minJ, comp909minVal, comp909minI, comp909minJ, comp2316minVal, comp2316minI, comp2316minJ);
    wire [11:0] comp2317minVal;
    wire [5:0] comp2317minI, comp2317minJ;
    Comparator comp2317(comp910minVal, comp910minI, comp910minJ, comp911minVal, comp911minI, comp911minJ, comp2317minVal, comp2317minI, comp2317minJ);
    wire [11:0] comp2318minVal;
    wire [5:0] comp2318minI, comp2318minJ;
    Comparator comp2318(comp912minVal, comp912minI, comp912minJ, comp913minVal, comp913minI, comp913minJ, comp2318minVal, comp2318minI, comp2318minJ);
    wire [11:0] comp2319minVal;
    wire [5:0] comp2319minI, comp2319minJ;
    Comparator comp2319(comp914minVal, comp914minI, comp914minJ, comp915minVal, comp915minI, comp915minJ, comp2319minVal, comp2319minI, comp2319minJ);
    wire [11:0] comp2320minVal;
    wire [5:0] comp2320minI, comp2320minJ;
    Comparator comp2320(comp916minVal, comp916minI, comp916minJ, comp917minVal, comp917minI, comp917minJ, comp2320minVal, comp2320minI, comp2320minJ);
    wire [11:0] comp2321minVal;
    wire [5:0] comp2321minI, comp2321minJ;
    Comparator comp2321(comp918minVal, comp918minI, comp918minJ, comp919minVal, comp919minI, comp919minJ, comp2321minVal, comp2321minI, comp2321minJ);
    wire [11:0] comp2322minVal;
    wire [5:0] comp2322minI, comp2322minJ;
    Comparator comp2322(comp920minVal, comp920minI, comp920minJ, comp921minVal, comp921minI, comp921minJ, comp2322minVal, comp2322minI, comp2322minJ);
    wire [11:0] comp2323minVal;
    wire [5:0] comp2323minI, comp2323minJ;
    Comparator comp2323(comp922minVal, comp922minI, comp922minJ, comp923minVal, comp923minI, comp923minJ, comp2323minVal, comp2323minI, comp2323minJ);
    wire [11:0] comp2324minVal;
    wire [5:0] comp2324minI, comp2324minJ;
    Comparator comp2324(comp924minVal, comp924minI, comp924minJ, comp925minVal, comp925minI, comp925minJ, comp2324minVal, comp2324minI, comp2324minJ);
    wire [11:0] comp2325minVal;
    wire [5:0] comp2325minI, comp2325minJ;
    Comparator comp2325(comp926minVal, comp926minI, comp926minJ, comp927minVal, comp927minI, comp927minJ, comp2325minVal, comp2325minI, comp2325minJ);
    wire [11:0] comp2326minVal;
    wire [5:0] comp2326minI, comp2326minJ;
    Comparator comp2326(comp928minVal, comp928minI, comp928minJ, comp929minVal, comp929minI, comp929minJ, comp2326minVal, comp2326minI, comp2326minJ);
    wire [11:0] comp2327minVal;
    wire [5:0] comp2327minI, comp2327minJ;
    Comparator comp2327(comp930minVal, comp930minI, comp930minJ, comp931minVal, comp931minI, comp931minJ, comp2327minVal, comp2327minI, comp2327minJ);
    wire [11:0] comp2328minVal;
    wire [5:0] comp2328minI, comp2328minJ;
    Comparator comp2328(comp932minVal, comp932minI, comp932minJ, comp933minVal, comp933minI, comp933minJ, comp2328minVal, comp2328minI, comp2328minJ);
    wire [11:0] comp2329minVal;
    wire [5:0] comp2329minI, comp2329minJ;
    Comparator comp2329(comp934minVal, comp934minI, comp934minJ, comp935minVal, comp935minI, comp935minJ, comp2329minVal, comp2329minI, comp2329minJ);
    wire [11:0] comp2330minVal;
    wire [5:0] comp2330minI, comp2330minJ;
    Comparator comp2330(comp936minVal, comp936minI, comp936minJ, comp937minVal, comp937minI, comp937minJ, comp2330minVal, comp2330minI, comp2330minJ);
    wire [11:0] comp2331minVal;
    wire [5:0] comp2331minI, comp2331minJ;
    Comparator comp2331(comp938minVal, comp938minI, comp938minJ, comp939minVal, comp939minI, comp939minJ, comp2331minVal, comp2331minI, comp2331minJ);
    wire [11:0] comp2332minVal;
    wire [5:0] comp2332minI, comp2332minJ;
    Comparator comp2332(comp940minVal, comp940minI, comp940minJ, comp941minVal, comp941minI, comp941minJ, comp2332minVal, comp2332minI, comp2332minJ);
    wire [11:0] comp2333minVal;
    wire [5:0] comp2333minI, comp2333minJ;
    Comparator comp2333(comp942minVal, comp942minI, comp942minJ, comp943minVal, comp943minI, comp943minJ, comp2333minVal, comp2333minI, comp2333minJ);
    wire [11:0] comp2334minVal;
    wire [5:0] comp2334minI, comp2334minJ;
    Comparator comp2334(comp944minVal, comp944minI, comp944minJ, comp945minVal, comp945minI, comp945minJ, comp2334minVal, comp2334minI, comp2334minJ);
    wire [11:0] comp2335minVal;
    wire [5:0] comp2335minI, comp2335minJ;
    Comparator comp2335(comp946minVal, comp946minI, comp946minJ, comp947minVal, comp947minI, comp947minJ, comp2335minVal, comp2335minI, comp2335minJ);
    wire [11:0] comp2336minVal;
    wire [5:0] comp2336minI, comp2336minJ;
    Comparator comp2336(comp948minVal, comp948minI, comp948minJ, comp949minVal, comp949minI, comp949minJ, comp2336minVal, comp2336minI, comp2336minJ);
    wire [11:0] comp2337minVal;
    wire [5:0] comp2337minI, comp2337minJ;
    Comparator comp2337(comp950minVal, comp950minI, comp950minJ, comp951minVal, comp951minI, comp951minJ, comp2337minVal, comp2337minI, comp2337minJ);
    wire [11:0] comp2338minVal;
    wire [5:0] comp2338minI, comp2338minJ;
    Comparator comp2338(comp952minVal, comp952minI, comp952minJ, comp953minVal, comp953minI, comp953minJ, comp2338minVal, comp2338minI, comp2338minJ);
    wire [11:0] comp2339minVal;
    wire [5:0] comp2339minI, comp2339minJ;
    Comparator comp2339(comp954minVal, comp954minI, comp954minJ, comp955minVal, comp955minI, comp955minJ, comp2339minVal, comp2339minI, comp2339minJ);
    wire [11:0] comp2340minVal;
    wire [5:0] comp2340minI, comp2340minJ;
    Comparator comp2340(comp956minVal, comp956minI, comp956minJ, comp957minVal, comp957minI, comp957minJ, comp2340minVal, comp2340minI, comp2340minJ);
    wire [11:0] comp2341minVal;
    wire [5:0] comp2341minI, comp2341minJ;
    Comparator comp2341(comp958minVal, comp958minI, comp958minJ, comp959minVal, comp959minI, comp959minJ, comp2341minVal, comp2341minI, comp2341minJ);
    wire [11:0] comp2342minVal;
    wire [5:0] comp2342minI, comp2342minJ;
    Comparator comp2342(comp960minVal, comp960minI, comp960minJ, comp961minVal, comp961minI, comp961minJ, comp2342minVal, comp2342minI, comp2342minJ);
    wire [11:0] comp2343minVal;
    wire [5:0] comp2343minI, comp2343minJ;
    Comparator comp2343(comp962minVal, comp962minI, comp962minJ, comp963minVal, comp963minI, comp963minJ, comp2343minVal, comp2343minI, comp2343minJ);
    wire [11:0] comp2344minVal;
    wire [5:0] comp2344minI, comp2344minJ;
    Comparator comp2344(comp964minVal, comp964minI, comp964minJ, comp965minVal, comp965minI, comp965minJ, comp2344minVal, comp2344minI, comp2344minJ);
    wire [11:0] comp2345minVal;
    wire [5:0] comp2345minI, comp2345minJ;
    Comparator comp2345(comp966minVal, comp966minI, comp966minJ, comp967minVal, comp967minI, comp967minJ, comp2345minVal, comp2345minI, comp2345minJ);
    wire [11:0] comp2346minVal;
    wire [5:0] comp2346minI, comp2346minJ;
    Comparator comp2346(comp968minVal, comp968minI, comp968minJ, comp969minVal, comp969minI, comp969minJ, comp2346minVal, comp2346minI, comp2346minJ);
    wire [11:0] comp2347minVal;
    wire [5:0] comp2347minI, comp2347minJ;
    Comparator comp2347(comp970minVal, comp970minI, comp970minJ, comp971minVal, comp971minI, comp971minJ, comp2347minVal, comp2347minI, comp2347minJ);
    wire [11:0] comp2348minVal;
    wire [5:0] comp2348minI, comp2348minJ;
    Comparator comp2348(comp972minVal, comp972minI, comp972minJ, comp973minVal, comp973minI, comp973minJ, comp2348minVal, comp2348minI, comp2348minJ);
    wire [11:0] comp2349minVal;
    wire [5:0] comp2349minI, comp2349minJ;
    Comparator comp2349(comp974minVal, comp974minI, comp974minJ, comp975minVal, comp975minI, comp975minJ, comp2349minVal, comp2349minI, comp2349minJ);
    wire [11:0] comp2350minVal;
    wire [5:0] comp2350minI, comp2350minJ;
    Comparator comp2350(comp976minVal, comp976minI, comp976minJ, comp977minVal, comp977minI, comp977minJ, comp2350minVal, comp2350minI, comp2350minJ);
    wire [11:0] comp2351minVal;
    wire [5:0] comp2351minI, comp2351minJ;
    Comparator comp2351(comp978minVal, comp978minI, comp978minJ, comp979minVal, comp979minI, comp979minJ, comp2351minVal, comp2351minI, comp2351minJ);
    wire [11:0] comp2352minVal;
    wire [5:0] comp2352minI, comp2352minJ;
    Comparator comp2352(comp980minVal, comp980minI, comp980minJ, comp981minVal, comp981minI, comp981minJ, comp2352minVal, comp2352minI, comp2352minJ);
    wire [11:0] comp2353minVal;
    wire [5:0] comp2353minI, comp2353minJ;
    Comparator comp2353(comp982minVal, comp982minI, comp982minJ, comp983minVal, comp983minI, comp983minJ, comp2353minVal, comp2353minI, comp2353minJ);
    wire [11:0] comp2354minVal;
    wire [5:0] comp2354minI, comp2354minJ;
    Comparator comp2354(comp984minVal, comp984minI, comp984minJ, comp985minVal, comp985minI, comp985minJ, comp2354minVal, comp2354minI, comp2354minJ);
    wire [11:0] comp2355minVal;
    wire [5:0] comp2355minI, comp2355minJ;
    Comparator comp2355(comp986minVal, comp986minI, comp986minJ, comp987minVal, comp987minI, comp987minJ, comp2355minVal, comp2355minI, comp2355minJ);
    wire [11:0] comp2356minVal;
    wire [5:0] comp2356minI, comp2356minJ;
    Comparator comp2356(comp988minVal, comp988minI, comp988minJ, comp989minVal, comp989minI, comp989minJ, comp2356minVal, comp2356minI, comp2356minJ);
    wire [11:0] comp2357minVal;
    wire [5:0] comp2357minI, comp2357minJ;
    Comparator comp2357(comp990minVal, comp990minI, comp990minJ, comp991minVal, comp991minI, comp991minJ, comp2357minVal, comp2357minI, comp2357minJ);
    wire [11:0] comp2358minVal;
    wire [5:0] comp2358minI, comp2358minJ;
    Comparator comp2358(comp992minVal, comp992minI, comp992minJ, comp993minVal, comp993minI, comp993minJ, comp2358minVal, comp2358minI, comp2358minJ);
    wire [11:0] comp2359minVal;
    wire [5:0] comp2359minI, comp2359minJ;
    Comparator comp2359(comp994minVal, comp994minI, comp994minJ, comp995minVal, comp995minI, comp995minJ, comp2359minVal, comp2359minI, comp2359minJ);
    wire [11:0] comp2360minVal;
    wire [5:0] comp2360minI, comp2360minJ;
    Comparator comp2360(comp996minVal, comp996minI, comp996minJ, comp997minVal, comp997minI, comp997minJ, comp2360minVal, comp2360minI, comp2360minJ);
    wire [11:0] comp2361minVal;
    wire [5:0] comp2361minI, comp2361minJ;
    Comparator comp2361(comp998minVal, comp998minI, comp998minJ, comp999minVal, comp999minI, comp999minJ, comp2361minVal, comp2361minI, comp2361minJ);
    wire [11:0] comp2362minVal;
    wire [5:0] comp2362minI, comp2362minJ;
    Comparator comp2362(comp1000minVal, comp1000minI, comp1000minJ, comp1001minVal, comp1001minI, comp1001minJ, comp2362minVal, comp2362minI, comp2362minJ);
    wire [11:0] comp2363minVal;
    wire [5:0] comp2363minI, comp2363minJ;
    Comparator comp2363(comp1002minVal, comp1002minI, comp1002minJ, comp1003minVal, comp1003minI, comp1003minJ, comp2363minVal, comp2363minI, comp2363minJ);
    wire [11:0] comp2364minVal;
    wire [5:0] comp2364minI, comp2364minJ;
    Comparator comp2364(comp1004minVal, comp1004minI, comp1004minJ, comp1005minVal, comp1005minI, comp1005minJ, comp2364minVal, comp2364minI, comp2364minJ);
    wire [11:0] comp2365minVal;
    wire [5:0] comp2365minI, comp2365minJ;
    Comparator comp2365(comp1006minVal, comp1006minI, comp1006minJ, comp1007minVal, comp1007minI, comp1007minJ, comp2365minVal, comp2365minI, comp2365minJ);
    wire [11:0] comp2366minVal;
    wire [5:0] comp2366minI, comp2366minJ;
    Comparator comp2366(comp1008minVal, comp1008minI, comp1008minJ, comp1009minVal, comp1009minI, comp1009minJ, comp2366minVal, comp2366minI, comp2366minJ);
    wire [11:0] comp2367minVal;
    wire [5:0] comp2367minI, comp2367minJ;
    Comparator comp2367(comp1010minVal, comp1010minI, comp1010minJ, comp1011minVal, comp1011minI, comp1011minJ, comp2367minVal, comp2367minI, comp2367minJ);
    wire [11:0] comp2368minVal;
    wire [5:0] comp2368minI, comp2368minJ;
    Comparator comp2368(comp1012minVal, comp1012minI, comp1012minJ, comp1013minVal, comp1013minI, comp1013minJ, comp2368minVal, comp2368minI, comp2368minJ);
    wire [11:0] comp2369minVal;
    wire [5:0] comp2369minI, comp2369minJ;
    Comparator comp2369(comp1014minVal, comp1014minI, comp1014minJ, comp1015minVal, comp1015minI, comp1015minJ, comp2369minVal, comp2369minI, comp2369minJ);
    wire [11:0] comp2370minVal;
    wire [5:0] comp2370minI, comp2370minJ;
    Comparator comp2370(comp1016minVal, comp1016minI, comp1016minJ, comp1017minVal, comp1017minI, comp1017minJ, comp2370minVal, comp2370minI, comp2370minJ);
    wire [11:0] comp2371minVal;
    wire [5:0] comp2371minI, comp2371minJ;
    Comparator comp2371(comp1018minVal, comp1018minI, comp1018minJ, comp1019minVal, comp1019minI, comp1019minJ, comp2371minVal, comp2371minI, comp2371minJ);
    wire [11:0] comp2372minVal;
    wire [5:0] comp2372minI, comp2372minJ;
    Comparator comp2372(comp1020minVal, comp1020minI, comp1020minJ, comp1021minVal, comp1021minI, comp1021minJ, comp2372minVal, comp2372minI, comp2372minJ);
    wire [11:0] comp2373minVal;
    wire [5:0] comp2373minI, comp2373minJ;
    Comparator comp2373(comp1022minVal, comp1022minI, comp1022minJ, comp1023minVal, comp1023minI, comp1023minJ, comp2373minVal, comp2373minI, comp2373minJ);
    wire [11:0] comp2374minVal;
    wire [5:0] comp2374minI, comp2374minJ;
    Comparator comp2374(comp1024minVal, comp1024minI, comp1024minJ, comp1025minVal, comp1025minI, comp1025minJ, comp2374minVal, comp2374minI, comp2374minJ);
    wire [11:0] comp2375minVal;
    wire [5:0] comp2375minI, comp2375minJ;
    Comparator comp2375(comp1026minVal, comp1026minI, comp1026minJ, comp1027minVal, comp1027minI, comp1027minJ, comp2375minVal, comp2375minI, comp2375minJ);
    wire [11:0] comp2376minVal;
    wire [5:0] comp2376minI, comp2376minJ;
    Comparator comp2376(comp1028minVal, comp1028minI, comp1028minJ, comp1029minVal, comp1029minI, comp1029minJ, comp2376minVal, comp2376minI, comp2376minJ);
    wire [11:0] comp2377minVal;
    wire [5:0] comp2377minI, comp2377minJ;
    Comparator comp2377(comp1030minVal, comp1030minI, comp1030minJ, comp1031minVal, comp1031minI, comp1031minJ, comp2377minVal, comp2377minI, comp2377minJ);
    wire [11:0] comp2378minVal;
    wire [5:0] comp2378minI, comp2378minJ;
    Comparator comp2378(comp1032minVal, comp1032minI, comp1032minJ, comp1033minVal, comp1033minI, comp1033minJ, comp2378minVal, comp2378minI, comp2378minJ);
    wire [11:0] comp2379minVal;
    wire [5:0] comp2379minI, comp2379minJ;
    Comparator comp2379(comp1034minVal, comp1034minI, comp1034minJ, comp1035minVal, comp1035minI, comp1035minJ, comp2379minVal, comp2379minI, comp2379minJ);
    wire [11:0] comp2380minVal;
    wire [5:0] comp2380minI, comp2380minJ;
    Comparator comp2380(comp1036minVal, comp1036minI, comp1036minJ, comp1037minVal, comp1037minI, comp1037minJ, comp2380minVal, comp2380minI, comp2380minJ);
    wire [11:0] comp2381minVal;
    wire [5:0] comp2381minI, comp2381minJ;
    Comparator comp2381(comp1038minVal, comp1038minI, comp1038minJ, comp1039minVal, comp1039minI, comp1039minJ, comp2381minVal, comp2381minI, comp2381minJ);
    wire [11:0] comp2382minVal;
    wire [5:0] comp2382minI, comp2382minJ;
    Comparator comp2382(comp1040minVal, comp1040minI, comp1040minJ, comp1041minVal, comp1041minI, comp1041minJ, comp2382minVal, comp2382minI, comp2382minJ);
    wire [11:0] comp2383minVal;
    wire [5:0] comp2383minI, comp2383minJ;
    Comparator comp2383(comp1042minVal, comp1042minI, comp1042minJ, comp1043minVal, comp1043minI, comp1043minJ, comp2383minVal, comp2383minI, comp2383minJ);
    wire [11:0] comp2384minVal;
    wire [5:0] comp2384minI, comp2384minJ;
    Comparator comp2384(comp1044minVal, comp1044minI, comp1044minJ, comp1045minVal, comp1045minI, comp1045minJ, comp2384minVal, comp2384minI, comp2384minJ);
    wire [11:0] comp2385minVal;
    wire [5:0] comp2385minI, comp2385minJ;
    Comparator comp2385(comp1046minVal, comp1046minI, comp1046minJ, comp1047minVal, comp1047minI, comp1047minJ, comp2385minVal, comp2385minI, comp2385minJ);
    wire [11:0] comp2386minVal;
    wire [5:0] comp2386minI, comp2386minJ;
    Comparator comp2386(comp1048minVal, comp1048minI, comp1048minJ, comp1049minVal, comp1049minI, comp1049minJ, comp2386minVal, comp2386minI, comp2386minJ);
    wire [11:0] comp2387minVal;
    wire [5:0] comp2387minI, comp2387minJ;
    Comparator comp2387(comp1050minVal, comp1050minI, comp1050minJ, comp1051minVal, comp1051minI, comp1051minJ, comp2387minVal, comp2387minI, comp2387minJ);
    wire [11:0] comp2388minVal;
    wire [5:0] comp2388minI, comp2388minJ;
    Comparator comp2388(comp1052minVal, comp1052minI, comp1052minJ, comp1053minVal, comp1053minI, comp1053minJ, comp2388minVal, comp2388minI, comp2388minJ);
    wire [11:0] comp2389minVal;
    wire [5:0] comp2389minI, comp2389minJ;
    Comparator comp2389(comp1054minVal, comp1054minI, comp1054minJ, comp1055minVal, comp1055minI, comp1055minJ, comp2389minVal, comp2389minI, comp2389minJ);
    wire [11:0] comp2390minVal;
    wire [5:0] comp2390minI, comp2390minJ;
    Comparator comp2390(comp1056minVal, comp1056minI, comp1056minJ, comp1057minVal, comp1057minI, comp1057minJ, comp2390minVal, comp2390minI, comp2390minJ);
    wire [11:0] comp2391minVal;
    wire [5:0] comp2391minI, comp2391minJ;
    Comparator comp2391(comp1058minVal, comp1058minI, comp1058minJ, comp1059minVal, comp1059minI, comp1059minJ, comp2391minVal, comp2391minI, comp2391minJ);
    wire [11:0] comp2392minVal;
    wire [5:0] comp2392minI, comp2392minJ;
    Comparator comp2392(comp1060minVal, comp1060minI, comp1060minJ, comp1061minVal, comp1061minI, comp1061minJ, comp2392minVal, comp2392minI, comp2392minJ);
    wire [11:0] comp2393minVal;
    wire [5:0] comp2393minI, comp2393minJ;
    Comparator comp2393(comp1062minVal, comp1062minI, comp1062minJ, comp1063minVal, comp1063minI, comp1063minJ, comp2393minVal, comp2393minI, comp2393minJ);
    wire [11:0] comp2394minVal;
    wire [5:0] comp2394minI, comp2394minJ;
    Comparator comp2394(comp1064minVal, comp1064minI, comp1064minJ, comp1065minVal, comp1065minI, comp1065minJ, comp2394minVal, comp2394minI, comp2394minJ);
    wire [11:0] comp2395minVal;
    wire [5:0] comp2395minI, comp2395minJ;
    Comparator comp2395(comp1066minVal, comp1066minI, comp1066minJ, comp1067minVal, comp1067minI, comp1067minJ, comp2395minVal, comp2395minI, comp2395minJ);
    wire [11:0] comp2396minVal;
    wire [5:0] comp2396minI, comp2396minJ;
    Comparator comp2396(comp1068minVal, comp1068minI, comp1068minJ, comp1069minVal, comp1069minI, comp1069minJ, comp2396minVal, comp2396minI, comp2396minJ);
    wire [11:0] comp2397minVal;
    wire [5:0] comp2397minI, comp2397minJ;
    Comparator comp2397(comp1070minVal, comp1070minI, comp1070minJ, comp1071minVal, comp1071minI, comp1071minJ, comp2397minVal, comp2397minI, comp2397minJ);
    wire [11:0] comp2398minVal;
    wire [5:0] comp2398minI, comp2398minJ;
    Comparator comp2398(comp1072minVal, comp1072minI, comp1072minJ, comp1073minVal, comp1073minI, comp1073minJ, comp2398minVal, comp2398minI, comp2398minJ);
    wire [11:0] comp2399minVal;
    wire [5:0] comp2399minI, comp2399minJ;
    Comparator comp2399(comp1074minVal, comp1074minI, comp1074minJ, comp1075minVal, comp1075minI, comp1075minJ, comp2399minVal, comp2399minI, comp2399minJ);
    wire [11:0] comp2400minVal;
    wire [5:0] comp2400minI, comp2400minJ;
    Comparator comp2400(comp1076minVal, comp1076minI, comp1076minJ, comp1077minVal, comp1077minI, comp1077minJ, comp2400minVal, comp2400minI, comp2400minJ);
    wire [11:0] comp2401minVal;
    wire [5:0] comp2401minI, comp2401minJ;
    Comparator comp2401(comp1078minVal, comp1078minI, comp1078minJ, comp1079minVal, comp1079minI, comp1079minJ, comp2401minVal, comp2401minI, comp2401minJ);
    wire [11:0] comp2402minVal;
    wire [5:0] comp2402minI, comp2402minJ;
    Comparator comp2402(comp1080minVal, comp1080minI, comp1080minJ, comp1081minVal, comp1081minI, comp1081minJ, comp2402minVal, comp2402minI, comp2402minJ);
    wire [11:0] comp2403minVal;
    wire [5:0] comp2403minI, comp2403minJ;
    Comparator comp2403(comp1082minVal, comp1082minI, comp1082minJ, comp1083minVal, comp1083minI, comp1083minJ, comp2403minVal, comp2403minI, comp2403minJ);
    wire [11:0] comp2404minVal;
    wire [5:0] comp2404minI, comp2404minJ;
    Comparator comp2404(comp1084minVal, comp1084minI, comp1084minJ, comp1085minVal, comp1085minI, comp1085minJ, comp2404minVal, comp2404minI, comp2404minJ);
    wire [11:0] comp2405minVal;
    wire [5:0] comp2405minI, comp2405minJ;
    Comparator comp2405(comp1086minVal, comp1086minI, comp1086minJ, comp1087minVal, comp1087minI, comp1087minJ, comp2405minVal, comp2405minI, comp2405minJ);
    wire [11:0] comp2406minVal;
    wire [5:0] comp2406minI, comp2406minJ;
    Comparator comp2406(comp1088minVal, comp1088minI, comp1088minJ, comp1089minVal, comp1089minI, comp1089minJ, comp2406minVal, comp2406minI, comp2406minJ);
    wire [11:0] comp2407minVal;
    wire [5:0] comp2407minI, comp2407minJ;
    Comparator comp2407(comp1090minVal, comp1090minI, comp1090minJ, comp1091minVal, comp1091minI, comp1091minJ, comp2407minVal, comp2407minI, comp2407minJ);
    wire [11:0] comp2408minVal;
    wire [5:0] comp2408minI, comp2408minJ;
    Comparator comp2408(comp1092minVal, comp1092minI, comp1092minJ, comp1093minVal, comp1093minI, comp1093minJ, comp2408minVal, comp2408minI, comp2408minJ);
    wire [11:0] comp2409minVal;
    wire [5:0] comp2409minI, comp2409minJ;
    Comparator comp2409(comp1094minVal, comp1094minI, comp1094minJ, comp1095minVal, comp1095minI, comp1095minJ, comp2409minVal, comp2409minI, comp2409minJ);
    wire [11:0] comp2410minVal;
    wire [5:0] comp2410minI, comp2410minJ;
    Comparator comp2410(comp1096minVal, comp1096minI, comp1096minJ, comp1097minVal, comp1097minI, comp1097minJ, comp2410minVal, comp2410minI, comp2410minJ);
    wire [11:0] comp2411minVal;
    wire [5:0] comp2411minI, comp2411minJ;
    Comparator comp2411(comp1098minVal, comp1098minI, comp1098minJ, comp1099minVal, comp1099minI, comp1099minJ, comp2411minVal, comp2411minI, comp2411minJ);
    wire [11:0] comp2412minVal;
    wire [5:0] comp2412minI, comp2412minJ;
    Comparator comp2412(comp1100minVal, comp1100minI, comp1100minJ, comp1101minVal, comp1101minI, comp1101minJ, comp2412minVal, comp2412minI, comp2412minJ);
    wire [11:0] comp2413minVal;
    wire [5:0] comp2413minI, comp2413minJ;
    Comparator comp2413(comp1102minVal, comp1102minI, comp1102minJ, comp1103minVal, comp1103minI, comp1103minJ, comp2413minVal, comp2413minI, comp2413minJ);
    wire [11:0] comp2414minVal;
    wire [5:0] comp2414minI, comp2414minJ;
    Comparator comp2414(comp1104minVal, comp1104minI, comp1104minJ, comp1105minVal, comp1105minI, comp1105minJ, comp2414minVal, comp2414minI, comp2414minJ);
    wire [11:0] comp2415minVal;
    wire [5:0] comp2415minI, comp2415minJ;
    Comparator comp2415(comp1106minVal, comp1106minI, comp1106minJ, comp1107minVal, comp1107minI, comp1107minJ, comp2415minVal, comp2415minI, comp2415minJ);
    wire [11:0] comp2416minVal;
    wire [5:0] comp2416minI, comp2416minJ;
    Comparator comp2416(comp1108minVal, comp1108minI, comp1108minJ, comp1109minVal, comp1109minI, comp1109minJ, comp2416minVal, comp2416minI, comp2416minJ);
    wire [11:0] comp2417minVal;
    wire [5:0] comp2417minI, comp2417minJ;
    Comparator comp2417(comp1110minVal, comp1110minI, comp1110minJ, comp1111minVal, comp1111minI, comp1111minJ, comp2417minVal, comp2417minI, comp2417minJ);
    wire [11:0] comp2418minVal;
    wire [5:0] comp2418minI, comp2418minJ;
    Comparator comp2418(comp1112minVal, comp1112minI, comp1112minJ, comp1113minVal, comp1113minI, comp1113minJ, comp2418minVal, comp2418minI, comp2418minJ);
    wire [11:0] comp2419minVal;
    wire [5:0] comp2419minI, comp2419minJ;
    Comparator comp2419(comp1114minVal, comp1114minI, comp1114minJ, comp1115minVal, comp1115minI, comp1115minJ, comp2419minVal, comp2419minI, comp2419minJ);
    wire [11:0] comp2420minVal;
    wire [5:0] comp2420minI, comp2420minJ;
    Comparator comp2420(comp1116minVal, comp1116minI, comp1116minJ, comp1117minVal, comp1117minI, comp1117minJ, comp2420minVal, comp2420minI, comp2420minJ);
    wire [11:0] comp2421minVal;
    wire [5:0] comp2421minI, comp2421minJ;
    Comparator comp2421(comp1118minVal, comp1118minI, comp1118minJ, comp1119minVal, comp1119minI, comp1119minJ, comp2421minVal, comp2421minI, comp2421minJ);
    wire [11:0] comp2422minVal;
    wire [5:0] comp2422minI, comp2422minJ;
    Comparator comp2422(comp1120minVal, comp1120minI, comp1120minJ, comp1121minVal, comp1121minI, comp1121minJ, comp2422minVal, comp2422minI, comp2422minJ);
    wire [11:0] comp2423minVal;
    wire [5:0] comp2423minI, comp2423minJ;
    Comparator comp2423(comp1122minVal, comp1122minI, comp1122minJ, comp1123minVal, comp1123minI, comp1123minJ, comp2423minVal, comp2423minI, comp2423minJ);
    wire [11:0] comp2424minVal;
    wire [5:0] comp2424minI, comp2424minJ;
    Comparator comp2424(comp1124minVal, comp1124minI, comp1124minJ, comp1125minVal, comp1125minI, comp1125minJ, comp2424minVal, comp2424minI, comp2424minJ);
    wire [11:0] comp2425minVal;
    wire [5:0] comp2425minI, comp2425minJ;
    Comparator comp2425(comp1126minVal, comp1126minI, comp1126minJ, comp1127minVal, comp1127minI, comp1127minJ, comp2425minVal, comp2425minI, comp2425minJ);
    wire [11:0] comp2426minVal;
    wire [5:0] comp2426minI, comp2426minJ;
    Comparator comp2426(comp1128minVal, comp1128minI, comp1128minJ, comp1129minVal, comp1129minI, comp1129minJ, comp2426minVal, comp2426minI, comp2426minJ);
    wire [11:0] comp2427minVal;
    wire [5:0] comp2427minI, comp2427minJ;
    Comparator comp2427(comp1130minVal, comp1130minI, comp1130minJ, comp1131minVal, comp1131minI, comp1131minJ, comp2427minVal, comp2427minI, comp2427minJ);
    wire [11:0] comp2428minVal;
    wire [5:0] comp2428minI, comp2428minJ;
    Comparator comp2428(comp1132minVal, comp1132minI, comp1132minJ, comp1133minVal, comp1133minI, comp1133minJ, comp2428minVal, comp2428minI, comp2428minJ);
    wire [11:0] comp2429minVal;
    wire [5:0] comp2429minI, comp2429minJ;
    Comparator comp2429(comp1134minVal, comp1134minI, comp1134minJ, comp1135minVal, comp1135minI, comp1135minJ, comp2429minVal, comp2429minI, comp2429minJ);
    wire [11:0] comp2430minVal;
    wire [5:0] comp2430minI, comp2430minJ;
    Comparator comp2430(comp1136minVal, comp1136minI, comp1136minJ, comp1137minVal, comp1137minI, comp1137minJ, comp2430minVal, comp2430minI, comp2430minJ);
    wire [11:0] comp2431minVal;
    wire [5:0] comp2431minI, comp2431minJ;
    Comparator comp2431(comp1138minVal, comp1138minI, comp1138minJ, comp1139minVal, comp1139minI, comp1139minJ, comp2431minVal, comp2431minI, comp2431minJ);
    wire [11:0] comp2432minVal;
    wire [5:0] comp2432minI, comp2432minJ;
    Comparator comp2432(comp1140minVal, comp1140minI, comp1140minJ, comp1141minVal, comp1141minI, comp1141minJ, comp2432minVal, comp2432minI, comp2432minJ);
    wire [11:0] comp2433minVal;
    wire [5:0] comp2433minI, comp2433minJ;
    Comparator comp2433(comp1142minVal, comp1142minI, comp1142minJ, comp1143minVal, comp1143minI, comp1143minJ, comp2433minVal, comp2433minI, comp2433minJ);
    wire [11:0] comp2434minVal;
    wire [5:0] comp2434minI, comp2434minJ;
    Comparator comp2434(comp1144minVal, comp1144minI, comp1144minJ, comp1145minVal, comp1145minI, comp1145minJ, comp2434minVal, comp2434minI, comp2434minJ);
    wire [11:0] comp2435minVal;
    wire [5:0] comp2435minI, comp2435minJ;
    Comparator comp2435(comp1146minVal, comp1146minI, comp1146minJ, comp1147minVal, comp1147minI, comp1147minJ, comp2435minVal, comp2435minI, comp2435minJ);
    wire [11:0] comp2436minVal;
    wire [5:0] comp2436minI, comp2436minJ;
    Comparator comp2436(comp1148minVal, comp1148minI, comp1148minJ, comp1149minVal, comp1149minI, comp1149minJ, comp2436minVal, comp2436minI, comp2436minJ);
    wire [11:0] comp2437minVal;
    wire [5:0] comp2437minI, comp2437minJ;
    Comparator comp2437(comp1150minVal, comp1150minI, comp1150minJ, comp1151minVal, comp1151minI, comp1151minJ, comp2437minVal, comp2437minI, comp2437minJ);
    wire [11:0] comp2438minVal;
    wire [5:0] comp2438minI, comp2438minJ;
    Comparator comp2438(comp1152minVal, comp1152minI, comp1152minJ, comp1153minVal, comp1153minI, comp1153minJ, comp2438minVal, comp2438minI, comp2438minJ);
    wire [11:0] comp2439minVal;
    wire [5:0] comp2439minI, comp2439minJ;
    Comparator comp2439(comp1154minVal, comp1154minI, comp1154minJ, comp1155minVal, comp1155minI, comp1155minJ, comp2439minVal, comp2439minI, comp2439minJ);
    wire [11:0] comp2440minVal;
    wire [5:0] comp2440minI, comp2440minJ;
    Comparator comp2440(comp1156minVal, comp1156minI, comp1156minJ, comp1157minVal, comp1157minI, comp1157minJ, comp2440minVal, comp2440minI, comp2440minJ);
    wire [11:0] comp2441minVal;
    wire [5:0] comp2441minI, comp2441minJ;
    Comparator comp2441(comp1158minVal, comp1158minI, comp1158minJ, comp1159minVal, comp1159minI, comp1159minJ, comp2441minVal, comp2441minI, comp2441minJ);
    wire [11:0] comp2442minVal;
    wire [5:0] comp2442minI, comp2442minJ;
    Comparator comp2442(comp1160minVal, comp1160minI, comp1160minJ, comp1161minVal, comp1161minI, comp1161minJ, comp2442minVal, comp2442minI, comp2442minJ);
    wire [11:0] comp2443minVal;
    wire [5:0] comp2443minI, comp2443minJ;
    Comparator comp2443(comp1162minVal, comp1162minI, comp1162minJ, comp1163minVal, comp1163minI, comp1163minJ, comp2443minVal, comp2443minI, comp2443minJ);
    wire [11:0] comp2444minVal;
    wire [5:0] comp2444minI, comp2444minJ;
    Comparator comp2444(comp1164minVal, comp1164minI, comp1164minJ, comp1165minVal, comp1165minI, comp1165minJ, comp2444minVal, comp2444minI, comp2444minJ);
    wire [11:0] comp2445minVal;
    wire [5:0] comp2445minI, comp2445minJ;
    Comparator comp2445(comp1166minVal, comp1166minI, comp1166minJ, comp1167minVal, comp1167minI, comp1167minJ, comp2445minVal, comp2445minI, comp2445minJ);
    wire [11:0] comp2446minVal;
    wire [5:0] comp2446minI, comp2446minJ;
    Comparator comp2446(comp1168minVal, comp1168minI, comp1168minJ, comp1169minVal, comp1169minI, comp1169minJ, comp2446minVal, comp2446minI, comp2446minJ);
    wire [11:0] comp2447minVal;
    wire [5:0] comp2447minI, comp2447minJ;
    Comparator comp2447(comp1170minVal, comp1170minI, comp1170minJ, comp1171minVal, comp1171minI, comp1171minJ, comp2447minVal, comp2447minI, comp2447minJ);
    wire [11:0] comp2448minVal;
    wire [5:0] comp2448minI, comp2448minJ;
    Comparator comp2448(comp1172minVal, comp1172minI, comp1172minJ, comp1173minVal, comp1173minI, comp1173minJ, comp2448minVal, comp2448minI, comp2448minJ);
    wire [11:0] comp2449minVal;
    wire [5:0] comp2449minI, comp2449minJ;
    Comparator comp2449(comp1174minVal, comp1174minI, comp1174minJ, comp1175minVal, comp1175minI, comp1175minJ, comp2449minVal, comp2449minI, comp2449minJ);
    wire [11:0] comp2450minVal;
    wire [5:0] comp2450minI, comp2450minJ;
    Comparator comp2450(comp1176minVal, comp1176minI, comp1176minJ, comp1177minVal, comp1177minI, comp1177minJ, comp2450minVal, comp2450minI, comp2450minJ);
    wire [11:0] comp2451minVal;
    wire [5:0] comp2451minI, comp2451minJ;
    Comparator comp2451(comp1178minVal, comp1178minI, comp1178minJ, comp1179minVal, comp1179minI, comp1179minJ, comp2451minVal, comp2451minI, comp2451minJ);
    wire [11:0] comp2452minVal;
    wire [5:0] comp2452minI, comp2452minJ;
    Comparator comp2452(comp1180minVal, comp1180minI, comp1180minJ, comp1181minVal, comp1181minI, comp1181minJ, comp2452minVal, comp2452minI, comp2452minJ);
    wire [11:0] comp2453minVal;
    wire [5:0] comp2453minI, comp2453minJ;
    Comparator comp2453(comp1182minVal, comp1182minI, comp1182minJ, comp1183minVal, comp1183minI, comp1183minJ, comp2453minVal, comp2453minI, comp2453minJ);
    wire [11:0] comp2454minVal;
    wire [5:0] comp2454minI, comp2454minJ;
    Comparator comp2454(comp1184minVal, comp1184minI, comp1184minJ, comp1185minVal, comp1185minI, comp1185minJ, comp2454minVal, comp2454minI, comp2454minJ);
    wire [11:0] comp2455minVal;
    wire [5:0] comp2455minI, comp2455minJ;
    Comparator comp2455(comp1186minVal, comp1186minI, comp1186minJ, comp1187minVal, comp1187minI, comp1187minJ, comp2455minVal, comp2455minI, comp2455minJ);
    wire [11:0] comp2456minVal;
    wire [5:0] comp2456minI, comp2456minJ;
    Comparator comp2456(comp1188minVal, comp1188minI, comp1188minJ, comp1189minVal, comp1189minI, comp1189minJ, comp2456minVal, comp2456minI, comp2456minJ);
    wire [11:0] comp2457minVal;
    wire [5:0] comp2457minI, comp2457minJ;
    Comparator comp2457(comp1190minVal, comp1190minI, comp1190minJ, comp1191minVal, comp1191minI, comp1191minJ, comp2457minVal, comp2457minI, comp2457minJ);
    wire [11:0] comp2458minVal;
    wire [5:0] comp2458minI, comp2458minJ;
    Comparator comp2458(comp1192minVal, comp1192minI, comp1192minJ, comp1193minVal, comp1193minI, comp1193minJ, comp2458minVal, comp2458minI, comp2458minJ);
    wire [11:0] comp2459minVal;
    wire [5:0] comp2459minI, comp2459minJ;
    Comparator comp2459(comp1194minVal, comp1194minI, comp1194minJ, comp1195minVal, comp1195minI, comp1195minJ, comp2459minVal, comp2459minI, comp2459minJ);
    wire [11:0] comp2460minVal;
    wire [5:0] comp2460minI, comp2460minJ;
    Comparator comp2460(comp1196minVal, comp1196minI, comp1196minJ, comp1197minVal, comp1197minI, comp1197minJ, comp2460minVal, comp2460minI, comp2460minJ);
    wire [11:0] comp2461minVal;
    wire [5:0] comp2461minI, comp2461minJ;
    Comparator comp2461(comp1198minVal, comp1198minI, comp1198minJ, comp1199minVal, comp1199minI, comp1199minJ, comp2461minVal, comp2461minI, comp2461minJ);
    wire [11:0] comp2462minVal;
    wire [5:0] comp2462minI, comp2462minJ;
    Comparator comp2462(comp1200minVal, comp1200minI, comp1200minJ, comp1201minVal, comp1201minI, comp1201minJ, comp2462minVal, comp2462minI, comp2462minJ);
    wire [11:0] comp2463minVal;
    wire [5:0] comp2463minI, comp2463minJ;
    Comparator comp2463(comp1202minVal, comp1202minI, comp1202minJ, comp1203minVal, comp1203minI, comp1203minJ, comp2463minVal, comp2463minI, comp2463minJ);
    wire [11:0] comp2464minVal;
    wire [5:0] comp2464minI, comp2464minJ;
    Comparator comp2464(comp1204minVal, comp1204minI, comp1204minJ, comp1205minVal, comp1205minI, comp1205minJ, comp2464minVal, comp2464minI, comp2464minJ);
    wire [11:0] comp2465minVal;
    wire [5:0] comp2465minI, comp2465minJ;
    Comparator comp2465(comp1206minVal, comp1206minI, comp1206minJ, comp1207minVal, comp1207minI, comp1207minJ, comp2465minVal, comp2465minI, comp2465minJ);
    wire [11:0] comp2466minVal;
    wire [5:0] comp2466minI, comp2466minJ;
    Comparator comp2466(comp1208minVal, comp1208minI, comp1208minJ, comp1209minVal, comp1209minI, comp1209minJ, comp2466minVal, comp2466minI, comp2466minJ);
    wire [11:0] comp2467minVal;
    wire [5:0] comp2467minI, comp2467minJ;
    Comparator comp2467(comp1210minVal, comp1210minI, comp1210minJ, comp1211minVal, comp1211minI, comp1211minJ, comp2467minVal, comp2467minI, comp2467minJ);
    wire [11:0] comp2468minVal;
    wire [5:0] comp2468minI, comp2468minJ;
    Comparator comp2468(comp1212minVal, comp1212minI, comp1212minJ, comp1213minVal, comp1213minI, comp1213minJ, comp2468minVal, comp2468minI, comp2468minJ);
    wire [11:0] comp2469minVal;
    wire [5:0] comp2469minI, comp2469minJ;
    Comparator comp2469(comp1214minVal, comp1214minI, comp1214minJ, comp1215minVal, comp1215minI, comp1215minJ, comp2469minVal, comp2469minI, comp2469minJ);
    wire [11:0] comp2470minVal;
    wire [5:0] comp2470minI, comp2470minJ;
    Comparator comp2470(comp1216minVal, comp1216minI, comp1216minJ, comp1217minVal, comp1217minI, comp1217minJ, comp2470minVal, comp2470minI, comp2470minJ);
    wire [11:0] comp2471minVal;
    wire [5:0] comp2471minI, comp2471minJ;
    Comparator comp2471(comp1218minVal, comp1218minI, comp1218minJ, comp1219minVal, comp1219minI, comp1219minJ, comp2471minVal, comp2471minI, comp2471minJ);
    wire [11:0] comp2472minVal;
    wire [5:0] comp2472minI, comp2472minJ;
    Comparator comp2472(comp1220minVal, comp1220minI, comp1220minJ, comp1221minVal, comp1221minI, comp1221minJ, comp2472minVal, comp2472minI, comp2472minJ);
    wire [11:0] comp2473minVal;
    wire [5:0] comp2473minI, comp2473minJ;
    Comparator comp2473(comp1222minVal, comp1222minI, comp1222minJ, comp1223minVal, comp1223minI, comp1223minJ, comp2473minVal, comp2473minI, comp2473minJ);
    wire [11:0] comp2474minVal;
    wire [5:0] comp2474minI, comp2474minJ;
    Comparator comp2474(comp1224minVal, comp1224minI, comp1224minJ, comp1225minVal, comp1225minI, comp1225minJ, comp2474minVal, comp2474minI, comp2474minJ);
    wire [11:0] comp2475minVal;
    wire [5:0] comp2475minI, comp2475minJ;
    Comparator comp2475(comp1226minVal, comp1226minI, comp1226minJ, comp1227minVal, comp1227minI, comp1227minJ, comp2475minVal, comp2475minI, comp2475minJ);
    wire [11:0] comp2476minVal;
    wire [5:0] comp2476minI, comp2476minJ;
    Comparator comp2476(comp1228minVal, comp1228minI, comp1228minJ, comp1229minVal, comp1229minI, comp1229minJ, comp2476minVal, comp2476minI, comp2476minJ);
    wire [11:0] comp2477minVal;
    wire [5:0] comp2477minI, comp2477minJ;
    Comparator comp2477(comp1230minVal, comp1230minI, comp1230minJ, comp1231minVal, comp1231minI, comp1231minJ, comp2477minVal, comp2477minI, comp2477minJ);
    wire [11:0] comp2478minVal;
    wire [5:0] comp2478minI, comp2478minJ;
    Comparator comp2478(comp1232minVal, comp1232minI, comp1232minJ, comp1233minVal, comp1233minI, comp1233minJ, comp2478minVal, comp2478minI, comp2478minJ);
    wire [11:0] comp2479minVal;
    wire [5:0] comp2479minI, comp2479minJ;
    Comparator comp2479(comp1234minVal, comp1234minI, comp1234minJ, comp1235minVal, comp1235minI, comp1235minJ, comp2479minVal, comp2479minI, comp2479minJ);
    wire [11:0] comp2480minVal;
    wire [5:0] comp2480minI, comp2480minJ;
    Comparator comp2480(comp1236minVal, comp1236minI, comp1236minJ, comp1237minVal, comp1237minI, comp1237minJ, comp2480minVal, comp2480minI, comp2480minJ);
    wire [11:0] comp2481minVal;
    wire [5:0] comp2481minI, comp2481minJ;
    Comparator comp2481(comp1238minVal, comp1238minI, comp1238minJ, comp1239minVal, comp1239minI, comp1239minJ, comp2481minVal, comp2481minI, comp2481minJ);
    wire [11:0] comp2482minVal;
    wire [5:0] comp2482minI, comp2482minJ;
    Comparator comp2482(comp1240minVal, comp1240minI, comp1240minJ, comp1241minVal, comp1241minI, comp1241minJ, comp2482minVal, comp2482minI, comp2482minJ);
    wire [11:0] comp2483minVal;
    wire [5:0] comp2483minI, comp2483minJ;
    Comparator comp2483(comp1242minVal, comp1242minI, comp1242minJ, comp1243minVal, comp1243minI, comp1243minJ, comp2483minVal, comp2483minI, comp2483minJ);
    wire [11:0] comp2484minVal;
    wire [5:0] comp2484minI, comp2484minJ;
    Comparator comp2484(comp1244minVal, comp1244minI, comp1244minJ, comp1245minVal, comp1245minI, comp1245minJ, comp2484minVal, comp2484minI, comp2484minJ);
    wire [11:0] comp2485minVal;
    wire [5:0] comp2485minI, comp2485minJ;
    Comparator comp2485(comp1246minVal, comp1246minI, comp1246minJ, comp1247minVal, comp1247minI, comp1247minJ, comp2485minVal, comp2485minI, comp2485minJ);
    wire [11:0] comp2486minVal;
    wire [5:0] comp2486minI, comp2486minJ;
    Comparator comp2486(comp1248minVal, comp1248minI, comp1248minJ, comp1249minVal, comp1249minI, comp1249minJ, comp2486minVal, comp2486minI, comp2486minJ);
    wire [11:0] comp2487minVal;
    wire [5:0] comp2487minI, comp2487minJ;
    Comparator comp2487(comp1250minVal, comp1250minI, comp1250minJ, comp1251minVal, comp1251minI, comp1251minJ, comp2487minVal, comp2487minI, comp2487minJ);
    wire [11:0] comp2488minVal;
    wire [5:0] comp2488minI, comp2488minJ;
    Comparator comp2488(comp1252minVal, comp1252minI, comp1252minJ, comp1253minVal, comp1253minI, comp1253minJ, comp2488minVal, comp2488minI, comp2488minJ);
    wire [11:0] comp2489minVal;
    wire [5:0] comp2489minI, comp2489minJ;
    Comparator comp2489(comp1254minVal, comp1254minI, comp1254minJ, comp1255minVal, comp1255minI, comp1255minJ, comp2489minVal, comp2489minI, comp2489minJ);
    wire [11:0] comp2490minVal;
    wire [5:0] comp2490minI, comp2490minJ;
    Comparator comp2490(comp1256minVal, comp1256minI, comp1256minJ, comp1257minVal, comp1257minI, comp1257minJ, comp2490minVal, comp2490minI, comp2490minJ);
    wire [11:0] comp2491minVal;
    wire [5:0] comp2491minI, comp2491minJ;
    Comparator comp2491(comp1258minVal, comp1258minI, comp1258minJ, comp1259minVal, comp1259minI, comp1259minJ, comp2491minVal, comp2491minI, comp2491minJ);
    wire [11:0] comp2492minVal;
    wire [5:0] comp2492minI, comp2492minJ;
    Comparator comp2492(comp1260minVal, comp1260minI, comp1260minJ, comp1261minVal, comp1261minI, comp1261minJ, comp2492minVal, comp2492minI, comp2492minJ);
    wire [11:0] comp2493minVal;
    wire [5:0] comp2493minI, comp2493minJ;
    Comparator comp2493(comp1262minVal, comp1262minI, comp1262minJ, comp1263minVal, comp1263minI, comp1263minJ, comp2493minVal, comp2493minI, comp2493minJ);
    wire [11:0] comp2494minVal;
    wire [5:0] comp2494minI, comp2494minJ;
    Comparator comp2494(comp1264minVal, comp1264minI, comp1264minJ, comp1265minVal, comp1265minI, comp1265minJ, comp2494minVal, comp2494minI, comp2494minJ);
    wire [11:0] comp2495minVal;
    wire [5:0] comp2495minI, comp2495minJ;
    Comparator comp2495(comp1266minVal, comp1266minI, comp1266minJ, comp1267minVal, comp1267minI, comp1267minJ, comp2495minVal, comp2495minI, comp2495minJ);
    wire [11:0] comp2496minVal;
    wire [5:0] comp2496minI, comp2496minJ;
    Comparator comp2496(comp1268minVal, comp1268minI, comp1268minJ, comp1269minVal, comp1269minI, comp1269minJ, comp2496minVal, comp2496minI, comp2496minJ);
    wire [11:0] comp2497minVal;
    wire [5:0] comp2497minI, comp2497minJ;
    Comparator comp2497(comp1270minVal, comp1270minI, comp1270minJ, comp1271minVal, comp1271minI, comp1271minJ, comp2497minVal, comp2497minI, comp2497minJ);
    wire [11:0] comp2498minVal;
    wire [5:0] comp2498minI, comp2498minJ;
    Comparator comp2498(comp1272minVal, comp1272minI, comp1272minJ, comp1273minVal, comp1273minI, comp1273minJ, comp2498minVal, comp2498minI, comp2498minJ);
    wire [11:0] comp2499minVal;
    wire [5:0] comp2499minI, comp2499minJ;
    Comparator comp2499(comp1274minVal, comp1274minI, comp1274minJ, comp1275minVal, comp1275minI, comp1275minJ, comp2499minVal, comp2499minI, comp2499minJ);
    wire [11:0] comp2500minVal;
    wire [5:0] comp2500minI, comp2500minJ;
    Comparator comp2500(comp1276minVal, comp1276minI, comp1276minJ, comp1277minVal, comp1277minI, comp1277minJ, comp2500minVal, comp2500minI, comp2500minJ);
    wire [11:0] comp2501minVal;
    wire [5:0] comp2501minI, comp2501minJ;
    Comparator comp2501(comp1278minVal, comp1278minI, comp1278minJ, comp1279minVal, comp1279minI, comp1279minJ, comp2501minVal, comp2501minI, comp2501minJ);
    wire [11:0] comp2502minVal;
    wire [5:0] comp2502minI, comp2502minJ;
    Comparator comp2502(comp1280minVal, comp1280minI, comp1280minJ, comp1281minVal, comp1281minI, comp1281minJ, comp2502minVal, comp2502minI, comp2502minJ);
    wire [11:0] comp2503minVal;
    wire [5:0] comp2503minI, comp2503minJ;
    Comparator comp2503(comp1282minVal, comp1282minI, comp1282minJ, comp1283minVal, comp1283minI, comp1283minJ, comp2503minVal, comp2503minI, comp2503minJ);
    wire [11:0] comp2504minVal;
    wire [5:0] comp2504minI, comp2504minJ;
    Comparator comp2504(comp1284minVal, comp1284minI, comp1284minJ, comp1285minVal, comp1285minI, comp1285minJ, comp2504minVal, comp2504minI, comp2504minJ);
    wire [11:0] comp2505minVal;
    wire [5:0] comp2505minI, comp2505minJ;
    Comparator comp2505(comp1286minVal, comp1286minI, comp1286minJ, comp1287minVal, comp1287minI, comp1287minJ, comp2505minVal, comp2505minI, comp2505minJ);
    wire [11:0] comp2506minVal;
    wire [5:0] comp2506minI, comp2506minJ;
    Comparator comp2506(comp1288minVal, comp1288minI, comp1288minJ, comp1289minVal, comp1289minI, comp1289minJ, comp2506minVal, comp2506minI, comp2506minJ);
    wire [11:0] comp2507minVal;
    wire [5:0] comp2507minI, comp2507minJ;
    Comparator comp2507(comp1290minVal, comp1290minI, comp1290minJ, comp1291minVal, comp1291minI, comp1291minJ, comp2507minVal, comp2507minI, comp2507minJ);
    wire [11:0] comp2508minVal;
    wire [5:0] comp2508minI, comp2508minJ;
    Comparator comp2508(comp1292minVal, comp1292minI, comp1292minJ, comp1293minVal, comp1293minI, comp1293minJ, comp2508minVal, comp2508minI, comp2508minJ);
    wire [11:0] comp2509minVal;
    wire [5:0] comp2509minI, comp2509minJ;
    Comparator comp2509(comp1294minVal, comp1294minI, comp1294minJ, comp1295minVal, comp1295minI, comp1295minJ, comp2509minVal, comp2509minI, comp2509minJ);
    wire [11:0] comp2510minVal;
    wire [5:0] comp2510minI, comp2510minJ;
    Comparator comp2510(comp1296minVal, comp1296minI, comp1296minJ, comp1297minVal, comp1297minI, comp1297minJ, comp2510minVal, comp2510minI, comp2510minJ);
    wire [11:0] comp2511minVal;
    wire [5:0] comp2511minI, comp2511minJ;
    Comparator comp2511(comp1298minVal, comp1298minI, comp1298minJ, comp1299minVal, comp1299minI, comp1299minJ, comp2511minVal, comp2511minI, comp2511minJ);
    wire [11:0] comp2512minVal;
    wire [5:0] comp2512minI, comp2512minJ;
    Comparator comp2512(comp1300minVal, comp1300minI, comp1300minJ, comp1301minVal, comp1301minI, comp1301minJ, comp2512minVal, comp2512minI, comp2512minJ);
    wire [11:0] comp2513minVal;
    wire [5:0] comp2513minI, comp2513minJ;
    Comparator comp2513(comp1302minVal, comp1302minI, comp1302minJ, comp1303minVal, comp1303minI, comp1303minJ, comp2513minVal, comp2513minI, comp2513minJ);
    wire [11:0] comp2514minVal;
    wire [5:0] comp2514minI, comp2514minJ;
    Comparator comp2514(comp1304minVal, comp1304minI, comp1304minJ, comp1305minVal, comp1305minI, comp1305minJ, comp2514minVal, comp2514minI, comp2514minJ);
    wire [11:0] comp2515minVal;
    wire [5:0] comp2515minI, comp2515minJ;
    Comparator comp2515(comp1306minVal, comp1306minI, comp1306minJ, comp1307minVal, comp1307minI, comp1307minJ, comp2515minVal, comp2515minI, comp2515minJ);
    wire [11:0] comp2516minVal;
    wire [5:0] comp2516minI, comp2516minJ;
    Comparator comp2516(comp1308minVal, comp1308minI, comp1308minJ, comp1309minVal, comp1309minI, comp1309minJ, comp2516minVal, comp2516minI, comp2516minJ);
    wire [11:0] comp2517minVal;
    wire [5:0] comp2517minI, comp2517minJ;
    Comparator comp2517(comp1310minVal, comp1310minI, comp1310minJ, comp1311minVal, comp1311minI, comp1311minJ, comp2517minVal, comp2517minI, comp2517minJ);
    wire [11:0] comp2518minVal;
    wire [5:0] comp2518minI, comp2518minJ;
    Comparator comp2518(comp1312minVal, comp1312minI, comp1312minJ, comp1313minVal, comp1313minI, comp1313minJ, comp2518minVal, comp2518minI, comp2518minJ);
    wire [11:0] comp2519minVal;
    wire [5:0] comp2519minI, comp2519minJ;
    Comparator comp2519(comp1314minVal, comp1314minI, comp1314minJ, comp1315minVal, comp1315minI, comp1315minJ, comp2519minVal, comp2519minI, comp2519minJ);
    wire [11:0] comp2520minVal;
    wire [5:0] comp2520minI, comp2520minJ;
    Comparator comp2520(comp1316minVal, comp1316minI, comp1316minJ, comp1317minVal, comp1317minI, comp1317minJ, comp2520minVal, comp2520minI, comp2520minJ);
    wire [11:0] comp2521minVal;
    wire [5:0] comp2521minI, comp2521minJ;
    Comparator comp2521(comp1318minVal, comp1318minI, comp1318minJ, comp1319minVal, comp1319minI, comp1319minJ, comp2521minVal, comp2521minI, comp2521minJ);
    wire [11:0] comp2522minVal;
    wire [5:0] comp2522minI, comp2522minJ;
    Comparator comp2522(comp1320minVal, comp1320minI, comp1320minJ, comp1321minVal, comp1321minI, comp1321minJ, comp2522minVal, comp2522minI, comp2522minJ);
    wire [11:0] comp2523minVal;
    wire [5:0] comp2523minI, comp2523minJ;
    Comparator comp2523(comp1322minVal, comp1322minI, comp1322minJ, comp1323minVal, comp1323minI, comp1323minJ, comp2523minVal, comp2523minI, comp2523minJ);
    wire [11:0] comp2524minVal;
    wire [5:0] comp2524minI, comp2524minJ;
    Comparator comp2524(comp1324minVal, comp1324minI, comp1324minJ, comp1325minVal, comp1325minI, comp1325minJ, comp2524minVal, comp2524minI, comp2524minJ);
    wire [11:0] comp2525minVal;
    wire [5:0] comp2525minI, comp2525minJ;
    Comparator comp2525(comp1326minVal, comp1326minI, comp1326minJ, comp1327minVal, comp1327minI, comp1327minJ, comp2525minVal, comp2525minI, comp2525minJ);
    wire [11:0] comp2526minVal;
    wire [5:0] comp2526minI, comp2526minJ;
    Comparator comp2526(comp1328minVal, comp1328minI, comp1328minJ, comp1329minVal, comp1329minI, comp1329minJ, comp2526minVal, comp2526minI, comp2526minJ);
    wire [11:0] comp2527minVal;
    wire [5:0] comp2527minI, comp2527minJ;
    Comparator comp2527(comp1330minVal, comp1330minI, comp1330minJ, comp1331minVal, comp1331minI, comp1331minJ, comp2527minVal, comp2527minI, comp2527minJ);
    wire [11:0] comp2528minVal;
    wire [5:0] comp2528minI, comp2528minJ;
    Comparator comp2528(comp1332minVal, comp1332minI, comp1332minJ, comp1333minVal, comp1333minI, comp1333minJ, comp2528minVal, comp2528minI, comp2528minJ);
    wire [11:0] comp2529minVal;
    wire [5:0] comp2529minI, comp2529minJ;
    Comparator comp2529(comp1334minVal, comp1334minI, comp1334minJ, comp1335minVal, comp1335minI, comp1335minJ, comp2529minVal, comp2529minI, comp2529minJ);
    wire [11:0] comp2530minVal;
    wire [5:0] comp2530minI, comp2530minJ;
    Comparator comp2530(comp1336minVal, comp1336minI, comp1336minJ, comp1337minVal, comp1337minI, comp1337minJ, comp2530minVal, comp2530minI, comp2530minJ);
    wire [11:0] comp2531minVal;
    wire [5:0] comp2531minI, comp2531minJ;
    Comparator comp2531(comp1338minVal, comp1338minI, comp1338minJ, comp1339minVal, comp1339minI, comp1339minJ, comp2531minVal, comp2531minI, comp2531minJ);
    wire [11:0] comp2532minVal;
    wire [5:0] comp2532minI, comp2532minJ;
    Comparator comp2532(comp1340minVal, comp1340minI, comp1340minJ, comp1341minVal, comp1341minI, comp1341minJ, comp2532minVal, comp2532minI, comp2532minJ);
    wire [11:0] comp2533minVal;
    wire [5:0] comp2533minI, comp2533minJ;
    Comparator comp2533(comp1342minVal, comp1342minI, comp1342minJ, comp1343minVal, comp1343minI, comp1343minJ, comp2533minVal, comp2533minI, comp2533minJ);
    wire [11:0] comp2534minVal;
    wire [5:0] comp2534minI, comp2534minJ;
    Comparator comp2534(comp1344minVal, comp1344minI, comp1344minJ, comp1345minVal, comp1345minI, comp1345minJ, comp2534minVal, comp2534minI, comp2534minJ);
    wire [11:0] comp2535minVal;
    wire [5:0] comp2535minI, comp2535minJ;
    Comparator comp2535(comp1346minVal, comp1346minI, comp1346minJ, comp1347minVal, comp1347minI, comp1347minJ, comp2535minVal, comp2535minI, comp2535minJ);
    wire [11:0] comp2536minVal;
    wire [5:0] comp2536minI, comp2536minJ;
    Comparator comp2536(comp1348minVal, comp1348minI, comp1348minJ, comp1349minVal, comp1349minI, comp1349minJ, comp2536minVal, comp2536minI, comp2536minJ);
    wire [11:0] comp2537minVal;
    wire [5:0] comp2537minI, comp2537minJ;
    Comparator comp2537(comp1350minVal, comp1350minI, comp1350minJ, comp1351minVal, comp1351minI, comp1351minJ, comp2537minVal, comp2537minI, comp2537minJ);
    wire [11:0] comp2538minVal;
    wire [5:0] comp2538minI, comp2538minJ;
    Comparator comp2538(comp1352minVal, comp1352minI, comp1352minJ, comp1353minVal, comp1353minI, comp1353minJ, comp2538minVal, comp2538minI, comp2538minJ);
    wire [11:0] comp2539minVal;
    wire [5:0] comp2539minI, comp2539minJ;
    Comparator comp2539(comp1354minVal, comp1354minI, comp1354minJ, comp1355minVal, comp1355minI, comp1355minJ, comp2539minVal, comp2539minI, comp2539minJ);
    wire [11:0] comp2540minVal;
    wire [5:0] comp2540minI, comp2540minJ;
    Comparator comp2540(comp1356minVal, comp1356minI, comp1356minJ, comp1357minVal, comp1357minI, comp1357minJ, comp2540minVal, comp2540minI, comp2540minJ);
    wire [11:0] comp2541minVal;
    wire [5:0] comp2541minI, comp2541minJ;
    Comparator comp2541(comp1358minVal, comp1358minI, comp1358minJ, comp1359minVal, comp1359minI, comp1359minJ, comp2541minVal, comp2541minI, comp2541minJ);
    wire [11:0] comp2542minVal;
    wire [5:0] comp2542minI, comp2542minJ;
    Comparator comp2542(comp1360minVal, comp1360minI, comp1360minJ, comp1361minVal, comp1361minI, comp1361minJ, comp2542minVal, comp2542minI, comp2542minJ);
    wire [11:0] comp2543minVal;
    wire [5:0] comp2543minI, comp2543minJ;
    Comparator comp2543(comp1362minVal, comp1362minI, comp1362minJ, comp1363minVal, comp1363minI, comp1363minJ, comp2543minVal, comp2543minI, comp2543minJ);
    wire [11:0] comp2544minVal;
    wire [5:0] comp2544minI, comp2544minJ;
    Comparator comp2544(comp1364minVal, comp1364minI, comp1364minJ, comp1365minVal, comp1365minI, comp1365minJ, comp2544minVal, comp2544minI, comp2544minJ);
    wire [11:0] comp2545minVal;
    wire [5:0] comp2545minI, comp2545minJ;
    Comparator comp2545(comp1366minVal, comp1366minI, comp1366minJ, comp1367minVal, comp1367minI, comp1367minJ, comp2545minVal, comp2545minI, comp2545minJ);
    wire [11:0] comp2546minVal;
    wire [5:0] comp2546minI, comp2546minJ;
    Comparator comp2546(comp1368minVal, comp1368minI, comp1368minJ, comp1369minVal, comp1369minI, comp1369minJ, comp2546minVal, comp2546minI, comp2546minJ);
    wire [11:0] comp2547minVal;
    wire [5:0] comp2547minI, comp2547minJ;
    Comparator comp2547(comp1370minVal, comp1370minI, comp1370minJ, comp1371minVal, comp1371minI, comp1371minJ, comp2547minVal, comp2547minI, comp2547minJ);
    wire [11:0] comp2548minVal;
    wire [5:0] comp2548minI, comp2548minJ;
    Comparator comp2548(comp1372minVal, comp1372minI, comp1372minJ, comp1373minVal, comp1373minI, comp1373minJ, comp2548minVal, comp2548minI, comp2548minJ);
    wire [11:0] comp2549minVal;
    wire [5:0] comp2549minI, comp2549minJ;
    Comparator comp2549(comp1374minVal, comp1374minI, comp1374minJ, comp1375minVal, comp1375minI, comp1375minJ, comp2549minVal, comp2549minI, comp2549minJ);
    wire [11:0] comp2550minVal;
    wire [5:0] comp2550minI, comp2550minJ;
    Comparator comp2550(comp1376minVal, comp1376minI, comp1376minJ, comp1377minVal, comp1377minI, comp1377minJ, comp2550minVal, comp2550minI, comp2550minJ);
    wire [11:0] comp2551minVal;
    wire [5:0] comp2551minI, comp2551minJ;
    Comparator comp2551(comp1378minVal, comp1378minI, comp1378minJ, comp1379minVal, comp1379minI, comp1379minJ, comp2551minVal, comp2551minI, comp2551minJ);
    wire [11:0] comp2552minVal;
    wire [5:0] comp2552minI, comp2552minJ;
    Comparator comp2552(comp1380minVal, comp1380minI, comp1380minJ, comp1381minVal, comp1381minI, comp1381minJ, comp2552minVal, comp2552minI, comp2552minJ);
    wire [11:0] comp2553minVal;
    wire [5:0] comp2553minI, comp2553minJ;
    Comparator comp2553(comp1382minVal, comp1382minI, comp1382minJ, comp1383minVal, comp1383minI, comp1383minJ, comp2553minVal, comp2553minI, comp2553minJ);
    wire [11:0] comp2554minVal;
    wire [5:0] comp2554minI, comp2554minJ;
    Comparator comp2554(comp1384minVal, comp1384minI, comp1384minJ, comp1385minVal, comp1385minI, comp1385minJ, comp2554minVal, comp2554minI, comp2554minJ);
    wire [11:0] comp2555minVal;
    wire [5:0] comp2555minI, comp2555minJ;
    Comparator comp2555(comp1386minVal, comp1386minI, comp1386minJ, comp1387minVal, comp1387minI, comp1387minJ, comp2555minVal, comp2555minI, comp2555minJ);
    wire [11:0] comp2556minVal;
    wire [5:0] comp2556minI, comp2556minJ;
    Comparator comp2556(comp1388minVal, comp1388minI, comp1388minJ, comp1389minVal, comp1389minI, comp1389minJ, comp2556minVal, comp2556minI, comp2556minJ);
    wire [11:0] comp2557minVal;
    wire [5:0] comp2557minI, comp2557minJ;
    Comparator comp2557(comp1390minVal, comp1390minI, comp1390minJ, comp1391minVal, comp1391minI, comp1391minJ, comp2557minVal, comp2557minI, comp2557minJ);
    wire [11:0] comp2558minVal;
    wire [5:0] comp2558minI, comp2558minJ;
    Comparator comp2558(comp1392minVal, comp1392minI, comp1392minJ, comp1393minVal, comp1393minI, comp1393minJ, comp2558minVal, comp2558minI, comp2558minJ);
    wire [11:0] comp2559minVal;
    wire [5:0] comp2559minI, comp2559minJ;
    Comparator comp2559(comp1394minVal, comp1394minI, comp1394minJ, comp1395minVal, comp1395minI, comp1395minJ, comp2559minVal, comp2559minI, comp2559minJ);
    wire [11:0] comp2560minVal;
    wire [5:0] comp2560minI, comp2560minJ;
    Comparator comp2560(comp1396minVal, comp1396minI, comp1396minJ, comp1397minVal, comp1397minI, comp1397minJ, comp2560minVal, comp2560minI, comp2560minJ);
    wire [11:0] comp2561minVal;
    wire [5:0] comp2561minI, comp2561minJ;
    Comparator comp2561(comp1398minVal, comp1398minI, comp1398minJ, comp1399minVal, comp1399minI, comp1399minJ, comp2561minVal, comp2561minI, comp2561minJ);
    wire [11:0] comp2562minVal;
    wire [5:0] comp2562minI, comp2562minJ;
    Comparator comp2562(comp1400minVal, comp1400minI, comp1400minJ, comp1401minVal, comp1401minI, comp1401minJ, comp2562minVal, comp2562minI, comp2562minJ);
    wire [11:0] comp2563minVal;
    wire [5:0] comp2563minI, comp2563minJ;
    Comparator comp2563(comp1402minVal, comp1402minI, comp1402minJ, comp1403minVal, comp1403minI, comp1403minJ, comp2563minVal, comp2563minI, comp2563minJ);
    wire [11:0] comp2564minVal;
    wire [5:0] comp2564minI, comp2564minJ;
    Comparator comp2564(comp1404minVal, comp1404minI, comp1404minJ, comp1405minVal, comp1405minI, comp1405minJ, comp2564minVal, comp2564minI, comp2564minJ);
    wire [11:0] comp2565minVal;
    wire [5:0] comp2565minI, comp2565minJ;
    Comparator comp2565(comp1406minVal, comp1406minI, comp1406minJ, comp1407minVal, comp1407minI, comp1407minJ, comp2565minVal, comp2565minI, comp2565minJ);
    wire [11:0] comp2566minVal;
    wire [5:0] comp2566minI, comp2566minJ;
    Comparator comp2566(comp1408minVal, comp1408minI, comp1408minJ, comp1409minVal, comp1409minI, comp1409minJ, comp2566minVal, comp2566minI, comp2566minJ);
    wire [11:0] comp2567minVal;
    wire [5:0] comp2567minI, comp2567minJ;
    Comparator comp2567(comp1410minVal, comp1410minI, comp1410minJ, comp1411minVal, comp1411minI, comp1411minJ, comp2567minVal, comp2567minI, comp2567minJ);
    wire [11:0] comp2568minVal;
    wire [5:0] comp2568minI, comp2568minJ;
    Comparator comp2568(comp1412minVal, comp1412minI, comp1412minJ, comp1413minVal, comp1413minI, comp1413minJ, comp2568minVal, comp2568minI, comp2568minJ);
    wire [11:0] comp2569minVal;
    wire [5:0] comp2569minI, comp2569minJ;
    Comparator comp2569(comp1414minVal, comp1414minI, comp1414minJ, comp1415minVal, comp1415minI, comp1415minJ, comp2569minVal, comp2569minI, comp2569minJ);
    wire [11:0] comp2570minVal;
    wire [5:0] comp2570minI, comp2570minJ;
    Comparator comp2570(comp1416minVal, comp1416minI, comp1416minJ, comp1417minVal, comp1417minI, comp1417minJ, comp2570minVal, comp2570minI, comp2570minJ);
    wire [11:0] comp2571minVal;
    wire [5:0] comp2571minI, comp2571minJ;
    Comparator comp2571(comp1418minVal, comp1418minI, comp1418minJ, comp1419minVal, comp1419minI, comp1419minJ, comp2571minVal, comp2571minI, comp2571minJ);
    wire [11:0] comp2572minVal;
    wire [5:0] comp2572minI, comp2572minJ;
    Comparator comp2572(comp1420minVal, comp1420minI, comp1420minJ, comp1421minVal, comp1421minI, comp1421minJ, comp2572minVal, comp2572minI, comp2572minJ);
    wire [11:0] comp2573minVal;
    wire [5:0] comp2573minI, comp2573minJ;
    Comparator comp2573(comp1422minVal, comp1422minI, comp1422minJ, comp1423minVal, comp1423minI, comp1423minJ, comp2573minVal, comp2573minI, comp2573minJ);
    wire [11:0] comp2574minVal;
    wire [5:0] comp2574minI, comp2574minJ;
    Comparator comp2574(comp1424minVal, comp1424minI, comp1424minJ, comp1425minVal, comp1425minI, comp1425minJ, comp2574minVal, comp2574minI, comp2574minJ);
    wire [11:0] comp2575minVal;
    wire [5:0] comp2575minI, comp2575minJ;
    Comparator comp2575(comp1426minVal, comp1426minI, comp1426minJ, comp1427minVal, comp1427minI, comp1427minJ, comp2575minVal, comp2575minI, comp2575minJ);
    wire [11:0] comp2576minVal;
    wire [5:0] comp2576minI, comp2576minJ;
    Comparator comp2576(comp1428minVal, comp1428minI, comp1428minJ, comp1429minVal, comp1429minI, comp1429minJ, comp2576minVal, comp2576minI, comp2576minJ);
    wire [11:0] comp2577minVal;
    wire [5:0] comp2577minI, comp2577minJ;
    Comparator comp2577(comp1430minVal, comp1430minI, comp1430minJ, comp1431minVal, comp1431minI, comp1431minJ, comp2577minVal, comp2577minI, comp2577minJ);
    wire [11:0] comp2578minVal;
    wire [5:0] comp2578minI, comp2578minJ;
    Comparator comp2578(comp1432minVal, comp1432minI, comp1432minJ, comp1433minVal, comp1433minI, comp1433minJ, comp2578minVal, comp2578minI, comp2578minJ);
    wire [11:0] comp2579minVal;
    wire [5:0] comp2579minI, comp2579minJ;
    Comparator comp2579(comp1434minVal, comp1434minI, comp1434minJ, comp1435minVal, comp1435minI, comp1435minJ, comp2579minVal, comp2579minI, comp2579minJ);
    wire [11:0] comp2580minVal;
    wire [5:0] comp2580minI, comp2580minJ;
    Comparator comp2580(comp1436minVal, comp1436minI, comp1436minJ, comp1437minVal, comp1437minI, comp1437minJ, comp2580minVal, comp2580minI, comp2580minJ);
    wire [11:0] comp2581minVal;
    wire [5:0] comp2581minI, comp2581minJ;
    Comparator comp2581(comp1438minVal, comp1438minI, comp1438minJ, comp1439minVal, comp1439minI, comp1439minJ, comp2581minVal, comp2581minI, comp2581minJ);
    wire [11:0] comp2582minVal;
    wire [5:0] comp2582minI, comp2582minJ;
    Comparator comp2582(comp1440minVal, comp1440minI, comp1440minJ, comp1441minVal, comp1441minI, comp1441minJ, comp2582minVal, comp2582minI, comp2582minJ);
    wire [11:0] comp2583minVal;
    wire [5:0] comp2583minI, comp2583minJ;
    Comparator comp2583(comp1442minVal, comp1442minI, comp1442minJ, comp1443minVal, comp1443minI, comp1443minJ, comp2583minVal, comp2583minI, comp2583minJ);
    wire [11:0] comp2584minVal;
    wire [5:0] comp2584minI, comp2584minJ;
    Comparator comp2584(comp1444minVal, comp1444minI, comp1444minJ, comp1445minVal, comp1445minI, comp1445minJ, comp2584minVal, comp2584minI, comp2584minJ);
    wire [11:0] comp2585minVal;
    wire [5:0] comp2585minI, comp2585minJ;
    Comparator comp2585(comp1446minVal, comp1446minI, comp1446minJ, comp1447minVal, comp1447minI, comp1447minJ, comp2585minVal, comp2585minI, comp2585minJ);
    wire [11:0] comp2586minVal;
    wire [5:0] comp2586minI, comp2586minJ;
    Comparator comp2586(comp1448minVal, comp1448minI, comp1448minJ, comp1449minVal, comp1449minI, comp1449minJ, comp2586minVal, comp2586minI, comp2586minJ);
    wire [11:0] comp2587minVal;
    wire [5:0] comp2587minI, comp2587minJ;
    Comparator comp2587(comp1450minVal, comp1450minI, comp1450minJ, comp1451minVal, comp1451minI, comp1451minJ, comp2587minVal, comp2587minI, comp2587minJ);
    wire [11:0] comp2588minVal;
    wire [5:0] comp2588minI, comp2588minJ;
    Comparator comp2588(comp1452minVal, comp1452minI, comp1452minJ, comp1453minVal, comp1453minI, comp1453minJ, comp2588minVal, comp2588minI, comp2588minJ);
    wire [11:0] comp2589minVal;
    wire [5:0] comp2589minI, comp2589minJ;
    Comparator comp2589(comp1454minVal, comp1454minI, comp1454minJ, comp1455minVal, comp1455minI, comp1455minJ, comp2589minVal, comp2589minI, comp2589minJ);
    wire [11:0] comp2590minVal;
    wire [5:0] comp2590minI, comp2590minJ;
    Comparator comp2590(comp1456minVal, comp1456minI, comp1456minJ, comp1457minVal, comp1457minI, comp1457minJ, comp2590minVal, comp2590minI, comp2590minJ);
    wire [11:0] comp2591minVal;
    wire [5:0] comp2591minI, comp2591minJ;
    Comparator comp2591(comp1458minVal, comp1458minI, comp1458minJ, comp1459minVal, comp1459minI, comp1459minJ, comp2591minVal, comp2591minI, comp2591minJ);
    wire [11:0] comp2592minVal;
    wire [5:0] comp2592minI, comp2592minJ;
    Comparator comp2592(comp1460minVal, comp1460minI, comp1460minJ, comp1461minVal, comp1461minI, comp1461minJ, comp2592minVal, comp2592minI, comp2592minJ);
    wire [11:0] comp2593minVal;
    wire [5:0] comp2593minI, comp2593minJ;
    Comparator comp2593(comp1462minVal, comp1462minI, comp1462minJ, comp1463minVal, comp1463minI, comp1463minJ, comp2593minVal, comp2593minI, comp2593minJ);
    wire [11:0] comp2594minVal;
    wire [5:0] comp2594minI, comp2594minJ;
    Comparator comp2594(comp1464minVal, comp1464minI, comp1464minJ, comp1465minVal, comp1465minI, comp1465minJ, comp2594minVal, comp2594minI, comp2594minJ);
    wire [11:0] comp2595minVal;
    wire [5:0] comp2595minI, comp2595minJ;
    Comparator comp2595(comp1466minVal, comp1466minI, comp1466minJ, comp1467minVal, comp1467minI, comp1467minJ, comp2595minVal, comp2595minI, comp2595minJ);
    wire [11:0] comp2596minVal;
    wire [5:0] comp2596minI, comp2596minJ;
    Comparator comp2596(comp1468minVal, comp1468minI, comp1468minJ, comp1469minVal, comp1469minI, comp1469minJ, comp2596minVal, comp2596minI, comp2596minJ);
    wire [11:0] comp2597minVal;
    wire [5:0] comp2597minI, comp2597minJ;
    Comparator comp2597(comp1470minVal, comp1470minI, comp1470minJ, comp1471minVal, comp1471minI, comp1471minJ, comp2597minVal, comp2597minI, comp2597minJ);
    wire [11:0] comp2598minVal;
    wire [5:0] comp2598minI, comp2598minJ;
    Comparator comp2598(comp1472minVal, comp1472minI, comp1472minJ, comp1473minVal, comp1473minI, comp1473minJ, comp2598minVal, comp2598minI, comp2598minJ);
    wire [11:0] comp2599minVal;
    wire [5:0] comp2599minI, comp2599minJ;
    Comparator comp2599(comp1474minVal, comp1474minI, comp1474minJ, comp1475minVal, comp1475minI, comp1475minJ, comp2599minVal, comp2599minI, comp2599minJ);
    wire [11:0] comp2600minVal;
    wire [5:0] comp2600minI, comp2600minJ;
    Comparator comp2600(comp1476minVal, comp1476minI, comp1476minJ, comp1477minVal, comp1477minI, comp1477minJ, comp2600minVal, comp2600minI, comp2600minJ);
    wire [11:0] comp2601minVal;
    wire [5:0] comp2601minI, comp2601minJ;
    Comparator comp2601(comp1478minVal, comp1478minI, comp1478minJ, comp1479minVal, comp1479minI, comp1479minJ, comp2601minVal, comp2601minI, comp2601minJ);
    wire [11:0] comp2602minVal;
    wire [5:0] comp2602minI, comp2602minJ;
    Comparator comp2602(comp1480minVal, comp1480minI, comp1480minJ, comp1481minVal, comp1481minI, comp1481minJ, comp2602minVal, comp2602minI, comp2602minJ);
    wire [11:0] comp2603minVal;
    wire [5:0] comp2603minI, comp2603minJ;
    Comparator comp2603(comp1482minVal, comp1482minI, comp1482minJ, comp1483minVal, comp1483minI, comp1483minJ, comp2603minVal, comp2603minI, comp2603minJ);
    wire [11:0] comp2604minVal;
    wire [5:0] comp2604minI, comp2604minJ;
    Comparator comp2604(comp1484minVal, comp1484minI, comp1484minJ, comp1485minVal, comp1485minI, comp1485minJ, comp2604minVal, comp2604minI, comp2604minJ);
    wire [11:0] comp2605minVal;
    wire [5:0] comp2605minI, comp2605minJ;
    Comparator comp2605(comp1486minVal, comp1486minI, comp1486minJ, comp1487minVal, comp1487minI, comp1487minJ, comp2605minVal, comp2605minI, comp2605minJ);
    wire [11:0] comp2606minVal;
    wire [5:0] comp2606minI, comp2606minJ;
    Comparator comp2606(comp1488minVal, comp1488minI, comp1488minJ, comp1489minVal, comp1489minI, comp1489minJ, comp2606minVal, comp2606minI, comp2606minJ);
    wire [11:0] comp2607minVal;
    wire [5:0] comp2607minI, comp2607minJ;
    Comparator comp2607(comp1490minVal, comp1490minI, comp1490minJ, comp1491minVal, comp1491minI, comp1491minJ, comp2607minVal, comp2607minI, comp2607minJ);
    wire [11:0] comp2608minVal;
    wire [5:0] comp2608minI, comp2608minJ;
    Comparator comp2608(comp1492minVal, comp1492minI, comp1492minJ, comp1493minVal, comp1493minI, comp1493minJ, comp2608minVal, comp2608minI, comp2608minJ);
    wire [11:0] comp2609minVal;
    wire [5:0] comp2609minI, comp2609minJ;
    Comparator comp2609(comp1494minVal, comp1494minI, comp1494minJ, comp1495minVal, comp1495minI, comp1495minJ, comp2609minVal, comp2609minI, comp2609minJ);
    wire [11:0] comp2610minVal;
    wire [5:0] comp2610minI, comp2610minJ;
    Comparator comp2610(comp1496minVal, comp1496minI, comp1496minJ, comp1497minVal, comp1497minI, comp1497minJ, comp2610minVal, comp2610minI, comp2610minJ);
    wire [11:0] comp2611minVal;
    wire [5:0] comp2611minI, comp2611minJ;
    Comparator comp2611(comp1498minVal, comp1498minI, comp1498minJ, comp1499minVal, comp1499minI, comp1499minJ, comp2611minVal, comp2611minI, comp2611minJ);
    wire [11:0] comp2612minVal;
    wire [5:0] comp2612minI, comp2612minJ;
    Comparator comp2612(comp1500minVal, comp1500minI, comp1500minJ, comp1501minVal, comp1501minI, comp1501minJ, comp2612minVal, comp2612minI, comp2612minJ);
    wire [11:0] comp2613minVal;
    wire [5:0] comp2613minI, comp2613minJ;
    Comparator comp2613(comp1502minVal, comp1502minI, comp1502minJ, comp1503minVal, comp1503minI, comp1503minJ, comp2613minVal, comp2613minI, comp2613minJ);
    wire [11:0] comp2614minVal;
    wire [5:0] comp2614minI, comp2614minJ;
    Comparator comp2614(comp1504minVal, comp1504minI, comp1504minJ, comp1505minVal, comp1505minI, comp1505minJ, comp2614minVal, comp2614minI, comp2614minJ);
    wire [11:0] comp2615minVal;
    wire [5:0] comp2615minI, comp2615minJ;
    Comparator comp2615(comp1506minVal, comp1506minI, comp1506minJ, comp1507minVal, comp1507minI, comp1507minJ, comp2615minVal, comp2615minI, comp2615minJ);
    wire [11:0] comp2616minVal;
    wire [5:0] comp2616minI, comp2616minJ;
    Comparator comp2616(comp1508minVal, comp1508minI, comp1508minJ, comp1509minVal, comp1509minI, comp1509minJ, comp2616minVal, comp2616minI, comp2616minJ);
    wire [11:0] comp2617minVal;
    wire [5:0] comp2617minI, comp2617minJ;
    Comparator comp2617(comp1510minVal, comp1510minI, comp1510minJ, comp1511minVal, comp1511minI, comp1511minJ, comp2617minVal, comp2617minI, comp2617minJ);
    wire [11:0] comp2618minVal;
    wire [5:0] comp2618minI, comp2618minJ;
    Comparator comp2618(comp1512minVal, comp1512minI, comp1512minJ, comp1513minVal, comp1513minI, comp1513minJ, comp2618minVal, comp2618minI, comp2618minJ);
    wire [11:0] comp2619minVal;
    wire [5:0] comp2619minI, comp2619minJ;
    Comparator comp2619(comp1514minVal, comp1514minI, comp1514minJ, comp1515minVal, comp1515minI, comp1515minJ, comp2619minVal, comp2619minI, comp2619minJ);
    wire [11:0] comp2620minVal;
    wire [5:0] comp2620minI, comp2620minJ;
    Comparator comp2620(comp1516minVal, comp1516minI, comp1516minJ, comp1517minVal, comp1517minI, comp1517minJ, comp2620minVal, comp2620minI, comp2620minJ);
    wire [11:0] comp2621minVal;
    wire [5:0] comp2621minI, comp2621minJ;
    Comparator comp2621(comp1518minVal, comp1518minI, comp1518minJ, comp1519minVal, comp1519minI, comp1519minJ, comp2621minVal, comp2621minI, comp2621minJ);
    wire [11:0] comp2622minVal;
    wire [5:0] comp2622minI, comp2622minJ;
    Comparator comp2622(comp1520minVal, comp1520minI, comp1520minJ, comp1521minVal, comp1521minI, comp1521minJ, comp2622minVal, comp2622minI, comp2622minJ);
    wire [11:0] comp2623minVal;
    wire [5:0] comp2623minI, comp2623minJ;
    Comparator comp2623(comp1522minVal, comp1522minI, comp1522minJ, comp1523minVal, comp1523minI, comp1523minJ, comp2623minVal, comp2623minI, comp2623minJ);
    wire [11:0] comp2624minVal;
    wire [5:0] comp2624minI, comp2624minJ;
    Comparator comp2624(comp1524minVal, comp1524minI, comp1524minJ, comp1525minVal, comp1525minI, comp1525minJ, comp2624minVal, comp2624minI, comp2624minJ);
    wire [11:0] comp2625minVal;
    wire [5:0] comp2625minI, comp2625minJ;
    Comparator comp2625(comp1526minVal, comp1526minI, comp1526minJ, comp1527minVal, comp1527minI, comp1527minJ, comp2625minVal, comp2625minI, comp2625minJ);
    wire [11:0] comp2626minVal;
    wire [5:0] comp2626minI, comp2626minJ;
    Comparator comp2626(comp1528minVal, comp1528minI, comp1528minJ, comp1529minVal, comp1529minI, comp1529minJ, comp2626minVal, comp2626minI, comp2626minJ);
    wire [11:0] comp2627minVal;
    wire [5:0] comp2627minI, comp2627minJ;
    Comparator comp2627(comp1530minVal, comp1530minI, comp1530minJ, comp1531minVal, comp1531minI, comp1531minJ, comp2627minVal, comp2627minI, comp2627minJ);
    wire [11:0] comp2628minVal;
    wire [5:0] comp2628minI, comp2628minJ;
    Comparator comp2628(comp1532minVal, comp1532minI, comp1532minJ, comp1533minVal, comp1533minI, comp1533minJ, comp2628minVal, comp2628minI, comp2628minJ);
    wire [11:0] comp2629minVal;
    wire [5:0] comp2629minI, comp2629minJ;
    Comparator comp2629(comp1534minVal, comp1534minI, comp1534minJ, comp1535minVal, comp1535minI, comp1535minJ, comp2629minVal, comp2629minI, comp2629minJ);
    wire [11:0] comp2630minVal;
    wire [5:0] comp2630minI, comp2630minJ;
    Comparator comp2630(comp1536minVal, comp1536minI, comp1536minJ, comp1537minVal, comp1537minI, comp1537minJ, comp2630minVal, comp2630minI, comp2630minJ);
    wire [11:0] comp2631minVal;
    wire [5:0] comp2631minI, comp2631minJ;
    Comparator comp2631(comp1538minVal, comp1538minI, comp1538minJ, comp1539minVal, comp1539minI, comp1539minJ, comp2631minVal, comp2631minI, comp2631minJ);
    wire [11:0] comp2632minVal;
    wire [5:0] comp2632minI, comp2632minJ;
    Comparator comp2632(comp1540minVal, comp1540minI, comp1540minJ, comp1541minVal, comp1541minI, comp1541minJ, comp2632minVal, comp2632minI, comp2632minJ);
    wire [11:0] comp2633minVal;
    wire [5:0] comp2633minI, comp2633minJ;
    Comparator comp2633(comp1542minVal, comp1542minI, comp1542minJ, comp1543minVal, comp1543minI, comp1543minJ, comp2633minVal, comp2633minI, comp2633minJ);
    wire [11:0] comp2634minVal;
    wire [5:0] comp2634minI, comp2634minJ;
    Comparator comp2634(comp1544minVal, comp1544minI, comp1544minJ, comp1545minVal, comp1545minI, comp1545minJ, comp2634minVal, comp2634minI, comp2634minJ);
    wire [11:0] comp2635minVal;
    wire [5:0] comp2635minI, comp2635minJ;
    Comparator comp2635(comp1546minVal, comp1546minI, comp1546minJ, comp1547minVal, comp1547minI, comp1547minJ, comp2635minVal, comp2635minI, comp2635minJ);
    wire [11:0] comp2636minVal;
    wire [5:0] comp2636minI, comp2636minJ;
    Comparator comp2636(comp1548minVal, comp1548minI, comp1548minJ, comp1549minVal, comp1549minI, comp1549minJ, comp2636minVal, comp2636minI, comp2636minJ);
    wire [11:0] comp2637minVal;
    wire [5:0] comp2637minI, comp2637minJ;
    Comparator comp2637(comp1550minVal, comp1550minI, comp1550minJ, comp1551minVal, comp1551minI, comp1551minJ, comp2637minVal, comp2637minI, comp2637minJ);
    wire [11:0] comp2638minVal;
    wire [5:0] comp2638minI, comp2638minJ;
    Comparator comp2638(comp1552minVal, comp1552minI, comp1552minJ, comp1553minVal, comp1553minI, comp1553minJ, comp2638minVal, comp2638minI, comp2638minJ);
    wire [11:0] comp2639minVal;
    wire [5:0] comp2639minI, comp2639minJ;
    Comparator comp2639(comp1554minVal, comp1554minI, comp1554minJ, comp1555minVal, comp1555minI, comp1555minJ, comp2639minVal, comp2639minI, comp2639minJ);
    wire [11:0] comp2640minVal;
    wire [5:0] comp2640minI, comp2640minJ;
    Comparator comp2640(comp1556minVal, comp1556minI, comp1556minJ, comp1557minVal, comp1557minI, comp1557minJ, comp2640minVal, comp2640minI, comp2640minJ);
    wire [11:0] comp2641minVal;
    wire [5:0] comp2641minI, comp2641minJ;
    Comparator comp2641(comp1558minVal, comp1558minI, comp1558minJ, comp1559minVal, comp1559minI, comp1559minJ, comp2641minVal, comp2641minI, comp2641minJ);
    wire [11:0] comp2642minVal;
    wire [5:0] comp2642minI, comp2642minJ;
    Comparator comp2642(comp1560minVal, comp1560minI, comp1560minJ, comp1561minVal, comp1561minI, comp1561minJ, comp2642minVal, comp2642minI, comp2642minJ);
    wire [11:0] comp2643minVal;
    wire [5:0] comp2643minI, comp2643minJ;
    Comparator comp2643(comp1562minVal, comp1562minI, comp1562minJ, comp1563minVal, comp1563minI, comp1563minJ, comp2643minVal, comp2643minI, comp2643minJ);
    wire [11:0] comp2644minVal;
    wire [5:0] comp2644minI, comp2644minJ;
    Comparator comp2644(comp1564minVal, comp1564minI, comp1564minJ, comp1565minVal, comp1565minI, comp1565minJ, comp2644minVal, comp2644minI, comp2644minJ);
    wire [11:0] comp2645minVal;
    wire [5:0] comp2645minI, comp2645minJ;
    Comparator comp2645(comp1566minVal, comp1566minI, comp1566minJ, comp1567minVal, comp1567minI, comp1567minJ, comp2645minVal, comp2645minI, comp2645minJ);
    wire [11:0] comp2646minVal;
    wire [5:0] comp2646minI, comp2646minJ;
    Comparator comp2646(comp1568minVal, comp1568minI, comp1568minJ, comp1569minVal, comp1569minI, comp1569minJ, comp2646minVal, comp2646minI, comp2646minJ);
    wire [11:0] comp2647minVal;
    wire [5:0] comp2647minI, comp2647minJ;
    Comparator comp2647(comp1570minVal, comp1570minI, comp1570minJ, comp1571minVal, comp1571minI, comp1571minJ, comp2647minVal, comp2647minI, comp2647minJ);
    wire [11:0] comp2648minVal;
    wire [5:0] comp2648minI, comp2648minJ;
    Comparator comp2648(comp1572minVal, comp1572minI, comp1572minJ, comp1573minVal, comp1573minI, comp1573minJ, comp2648minVal, comp2648minI, comp2648minJ);
    wire [11:0] comp2649minVal;
    wire [5:0] comp2649minI, comp2649minJ;
    Comparator comp2649(comp1574minVal, comp1574minI, comp1574minJ, comp1575minVal, comp1575minI, comp1575minJ, comp2649minVal, comp2649minI, comp2649minJ);
    wire [11:0] comp2650minVal;
    wire [5:0] comp2650minI, comp2650minJ;
    Comparator comp2650(comp1576minVal, comp1576minI, comp1576minJ, comp1577minVal, comp1577minI, comp1577minJ, comp2650minVal, comp2650minI, comp2650minJ);
    wire [11:0] comp2651minVal;
    wire [5:0] comp2651minI, comp2651minJ;
    Comparator comp2651(comp1578minVal, comp1578minI, comp1578minJ, comp1579minVal, comp1579minI, comp1579minJ, comp2651minVal, comp2651minI, comp2651minJ);
    wire [11:0] comp2652minVal;
    wire [5:0] comp2652minI, comp2652minJ;
    Comparator comp2652(comp1580minVal, comp1580minI, comp1580minJ, comp1581minVal, comp1581minI, comp1581minJ, comp2652minVal, comp2652minI, comp2652minJ);
    wire [11:0] comp2653minVal;
    wire [5:0] comp2653minI, comp2653minJ;
    Comparator comp2653(comp1582minVal, comp1582minI, comp1582minJ, comp1583minVal, comp1583minI, comp1583minJ, comp2653minVal, comp2653minI, comp2653minJ);
    wire [11:0] comp2654minVal;
    wire [5:0] comp2654minI, comp2654minJ;
    Comparator comp2654(comp1584minVal, comp1584minI, comp1584minJ, comp1585minVal, comp1585minI, comp1585minJ, comp2654minVal, comp2654minI, comp2654minJ);
    wire [11:0] comp2655minVal;
    wire [5:0] comp2655minI, comp2655minJ;
    Comparator comp2655(comp1586minVal, comp1586minI, comp1586minJ, comp1587minVal, comp1587minI, comp1587minJ, comp2655minVal, comp2655minI, comp2655minJ);
    wire [11:0] comp2656minVal;
    wire [5:0] comp2656minI, comp2656minJ;
    Comparator comp2656(comp1588minVal, comp1588minI, comp1588minJ, comp1589minVal, comp1589minI, comp1589minJ, comp2656minVal, comp2656minI, comp2656minJ);
    wire [11:0] comp2657minVal;
    wire [5:0] comp2657minI, comp2657minJ;
    Comparator comp2657(comp1590minVal, comp1590minI, comp1590minJ, comp1591minVal, comp1591minI, comp1591minJ, comp2657minVal, comp2657minI, comp2657minJ);
    wire [11:0] comp2658minVal;
    wire [5:0] comp2658minI, comp2658minJ;
    Comparator comp2658(comp1592minVal, comp1592minI, comp1592minJ, comp1593minVal, comp1593minI, comp1593minJ, comp2658minVal, comp2658minI, comp2658minJ);
    wire [11:0] comp2659minVal;
    wire [5:0] comp2659minI, comp2659minJ;
    Comparator comp2659(comp1594minVal, comp1594minI, comp1594minJ, comp1595minVal, comp1595minI, comp1595minJ, comp2659minVal, comp2659minI, comp2659minJ);
    wire [11:0] comp2660minVal;
    wire [5:0] comp2660minI, comp2660minJ;
    Comparator comp2660(comp1596minVal, comp1596minI, comp1596minJ, comp1597minVal, comp1597minI, comp1597minJ, comp2660minVal, comp2660minI, comp2660minJ);
    wire [11:0] comp2661minVal;
    wire [5:0] comp2661minI, comp2661minJ;
    Comparator comp2661(comp1598minVal, comp1598minI, comp1598minJ, comp1599minVal, comp1599minI, comp1599minJ, comp2661minVal, comp2661minI, comp2661minJ);
    wire [11:0] comp2662minVal;
    wire [5:0] comp2662minI, comp2662minJ;
    Comparator comp2662(comp1600minVal, comp1600minI, comp1600minJ, comp1601minVal, comp1601minI, comp1601minJ, comp2662minVal, comp2662minI, comp2662minJ);
    wire [11:0] comp2663minVal;
    wire [5:0] comp2663minI, comp2663minJ;
    Comparator comp2663(comp1602minVal, comp1602minI, comp1602minJ, comp1603minVal, comp1603minI, comp1603minJ, comp2663minVal, comp2663minI, comp2663minJ);
    wire [11:0] comp2664minVal;
    wire [5:0] comp2664minI, comp2664minJ;
    Comparator comp2664(comp1604minVal, comp1604minI, comp1604minJ, comp1605minVal, comp1605minI, comp1605minJ, comp2664minVal, comp2664minI, comp2664minJ);
    wire [11:0] comp2665minVal;
    wire [5:0] comp2665minI, comp2665minJ;
    Comparator comp2665(comp1606minVal, comp1606minI, comp1606minJ, comp1607minVal, comp1607minI, comp1607minJ, comp2665minVal, comp2665minI, comp2665minJ);
    wire [11:0] comp2666minVal;
    wire [5:0] comp2666minI, comp2666minJ;
    Comparator comp2666(comp1608minVal, comp1608minI, comp1608minJ, comp1609minVal, comp1609minI, comp1609minJ, comp2666minVal, comp2666minI, comp2666minJ);
    wire [11:0] comp2667minVal;
    wire [5:0] comp2667minI, comp2667minJ;
    Comparator comp2667(comp1610minVal, comp1610minI, comp1610minJ, comp1611minVal, comp1611minI, comp1611minJ, comp2667minVal, comp2667minI, comp2667minJ);
    wire [11:0] comp2668minVal;
    wire [5:0] comp2668minI, comp2668minJ;
    Comparator comp2668(comp1612minVal, comp1612minI, comp1612minJ, comp1613minVal, comp1613minI, comp1613minJ, comp2668minVal, comp2668minI, comp2668minJ);
    wire [11:0] comp2669minVal;
    wire [5:0] comp2669minI, comp2669minJ;
    Comparator comp2669(comp1614minVal, comp1614minI, comp1614minJ, comp1615minVal, comp1615minI, comp1615minJ, comp2669minVal, comp2669minI, comp2669minJ);
    wire [11:0] comp2670minVal;
    wire [5:0] comp2670minI, comp2670minJ;
    Comparator comp2670(comp1616minVal, comp1616minI, comp1616minJ, comp1617minVal, comp1617minI, comp1617minJ, comp2670minVal, comp2670minI, comp2670minJ);
    wire [11:0] comp2671minVal;
    wire [5:0] comp2671minI, comp2671minJ;
    Comparator comp2671(comp1618minVal, comp1618minI, comp1618minJ, comp1619minVal, comp1619minI, comp1619minJ, comp2671minVal, comp2671minI, comp2671minJ);
    wire [11:0] comp2672minVal;
    wire [5:0] comp2672minI, comp2672minJ;
    Comparator comp2672(comp1620minVal, comp1620minI, comp1620minJ, comp1621minVal, comp1621minI, comp1621minJ, comp2672minVal, comp2672minI, comp2672minJ);
    wire [11:0] comp2673minVal;
    wire [5:0] comp2673minI, comp2673minJ;
    Comparator comp2673(comp1622minVal, comp1622minI, comp1622minJ, comp1623minVal, comp1623minI, comp1623minJ, comp2673minVal, comp2673minI, comp2673minJ);
    wire [11:0] comp2674minVal;
    wire [5:0] comp2674minI, comp2674minJ;
    Comparator comp2674(comp1624minVal, comp1624minI, comp1624minJ, comp1625minVal, comp1625minI, comp1625minJ, comp2674minVal, comp2674minI, comp2674minJ);
    wire [11:0] comp2675minVal;
    wire [5:0] comp2675minI, comp2675minJ;
    Comparator comp2675(comp1626minVal, comp1626minI, comp1626minJ, comp1627minVal, comp1627minI, comp1627minJ, comp2675minVal, comp2675minI, comp2675minJ);
    wire [11:0] comp2676minVal;
    wire [5:0] comp2676minI, comp2676minJ;
    Comparator comp2676(comp1628minVal, comp1628minI, comp1628minJ, comp1629minVal, comp1629minI, comp1629minJ, comp2676minVal, comp2676minI, comp2676minJ);
    wire [11:0] comp2677minVal;
    wire [5:0] comp2677minI, comp2677minJ;
    Comparator comp2677(comp1630minVal, comp1630minI, comp1630minJ, comp1631minVal, comp1631minI, comp1631minJ, comp2677minVal, comp2677minI, comp2677minJ);
    wire [11:0] comp2678minVal;
    wire [5:0] comp2678minI, comp2678minJ;
    Comparator comp2678(comp1632minVal, comp1632minI, comp1632minJ, comp1633minVal, comp1633minI, comp1633minJ, comp2678minVal, comp2678minI, comp2678minJ);
    wire [11:0] comp2679minVal;
    wire [5:0] comp2679minI, comp2679minJ;
    Comparator comp2679(comp1634minVal, comp1634minI, comp1634minJ, comp1635minVal, comp1635minI, comp1635minJ, comp2679minVal, comp2679minI, comp2679minJ);
    wire [11:0] comp2680minVal;
    wire [5:0] comp2680minI, comp2680minJ;
    Comparator comp2680(comp1636minVal, comp1636minI, comp1636minJ, comp1637minVal, comp1637minI, comp1637minJ, comp2680minVal, comp2680minI, comp2680minJ);
    wire [11:0] comp2681minVal;
    wire [5:0] comp2681minI, comp2681minJ;
    Comparator comp2681(comp1638minVal, comp1638minI, comp1638minJ, comp1639minVal, comp1639minI, comp1639minJ, comp2681minVal, comp2681minI, comp2681minJ);
    wire [11:0] comp2682minVal;
    wire [5:0] comp2682minI, comp2682minJ;
    Comparator comp2682(comp1640minVal, comp1640minI, comp1640minJ, comp1641minVal, comp1641minI, comp1641minJ, comp2682minVal, comp2682minI, comp2682minJ);
    wire [11:0] comp2683minVal;
    wire [5:0] comp2683minI, comp2683minJ;
    Comparator comp2683(comp1642minVal, comp1642minI, comp1642minJ, comp1643minVal, comp1643minI, comp1643minJ, comp2683minVal, comp2683minI, comp2683minJ);
    wire [11:0] comp2684minVal;
    wire [5:0] comp2684minI, comp2684minJ;
    Comparator comp2684(comp1644minVal, comp1644minI, comp1644minJ, comp1645minVal, comp1645minI, comp1645minJ, comp2684minVal, comp2684minI, comp2684minJ);
    wire [11:0] comp2685minVal;
    wire [5:0] comp2685minI, comp2685minJ;
    Comparator comp2685(comp1646minVal, comp1646minI, comp1646minJ, comp1647minVal, comp1647minI, comp1647minJ, comp2685minVal, comp2685minI, comp2685minJ);
    wire [11:0] comp2686minVal;
    wire [5:0] comp2686minI, comp2686minJ;
    Comparator comp2686(comp1648minVal, comp1648minI, comp1648minJ, comp1649minVal, comp1649minI, comp1649minJ, comp2686minVal, comp2686minI, comp2686minJ);
    wire [11:0] comp2687minVal;
    wire [5:0] comp2687minI, comp2687minJ;
    Comparator comp2687(comp1650minVal, comp1650minI, comp1650minJ, comp1651minVal, comp1651minI, comp1651minJ, comp2687minVal, comp2687minI, comp2687minJ);
    wire [11:0] comp2688minVal;
    wire [5:0] comp2688minI, comp2688minJ;
    Comparator comp2688(comp1652minVal, comp1652minI, comp1652minJ, comp1653minVal, comp1653minI, comp1653minJ, comp2688minVal, comp2688minI, comp2688minJ);
    wire [11:0] comp2689minVal;
    wire [5:0] comp2689minI, comp2689minJ;
    Comparator comp2689(comp1654minVal, comp1654minI, comp1654minJ, comp1655minVal, comp1655minI, comp1655minJ, comp2689minVal, comp2689minI, comp2689minJ);
    wire [11:0] comp2690minVal;
    wire [5:0] comp2690minI, comp2690minJ;
    Comparator comp2690(comp1656minVal, comp1656minI, comp1656minJ, comp1657minVal, comp1657minI, comp1657minJ, comp2690minVal, comp2690minI, comp2690minJ);
    wire [11:0] comp2691minVal;
    wire [5:0] comp2691minI, comp2691minJ;
    Comparator comp2691(comp1658minVal, comp1658minI, comp1658minJ, comp1659minVal, comp1659minI, comp1659minJ, comp2691minVal, comp2691minI, comp2691minJ);
    wire [11:0] comp2692minVal;
    wire [5:0] comp2692minI, comp2692minJ;
    Comparator comp2692(comp1660minVal, comp1660minI, comp1660minJ, comp1661minVal, comp1661minI, comp1661minJ, comp2692minVal, comp2692minI, comp2692minJ);
    wire [11:0] comp2693minVal;
    wire [5:0] comp2693minI, comp2693minJ;
    Comparator comp2693(comp1662minVal, comp1662minI, comp1662minJ, comp1663minVal, comp1663minI, comp1663minJ, comp2693minVal, comp2693minI, comp2693minJ);
    wire [11:0] comp2694minVal;
    wire [5:0] comp2694minI, comp2694minJ;
    Comparator comp2694(comp1664minVal, comp1664minI, comp1664minJ, comp1665minVal, comp1665minI, comp1665minJ, comp2694minVal, comp2694minI, comp2694minJ);
    wire [11:0] comp2695minVal;
    wire [5:0] comp2695minI, comp2695minJ;
    Comparator comp2695(comp1666minVal, comp1666minI, comp1666minJ, comp1667minVal, comp1667minI, comp1667minJ, comp2695minVal, comp2695minI, comp2695minJ);
    wire [11:0] comp2696minVal;
    wire [5:0] comp2696minI, comp2696minJ;
    Comparator comp2696(comp1668minVal, comp1668minI, comp1668minJ, comp1669minVal, comp1669minI, comp1669minJ, comp2696minVal, comp2696minI, comp2696minJ);
    wire [11:0] comp2697minVal;
    wire [5:0] comp2697minI, comp2697minJ;
    Comparator comp2697(comp1670minVal, comp1670minI, comp1670minJ, comp1671minVal, comp1671minI, comp1671minJ, comp2697minVal, comp2697minI, comp2697minJ);
    wire [11:0] comp2698minVal;
    wire [5:0] comp2698minI, comp2698minJ;
    Comparator comp2698(comp1672minVal, comp1672minI, comp1672minJ, comp1673minVal, comp1673minI, comp1673minJ, comp2698minVal, comp2698minI, comp2698minJ);
    wire [11:0] comp2699minVal;
    wire [5:0] comp2699minI, comp2699minJ;
    Comparator comp2699(comp1674minVal, comp1674minI, comp1674minJ, comp1675minVal, comp1675minI, comp1675minJ, comp2699minVal, comp2699minI, comp2699minJ);
    wire [11:0] comp2700minVal;
    wire [5:0] comp2700minI, comp2700minJ;
    Comparator comp2700(comp1676minVal, comp1676minI, comp1676minJ, comp1677minVal, comp1677minI, comp1677minJ, comp2700minVal, comp2700minI, comp2700minJ);
    wire [11:0] comp2701minVal;
    wire [5:0] comp2701minI, comp2701minJ;
    Comparator comp2701(comp1678minVal, comp1678minI, comp1678minJ, comp1679minVal, comp1679minI, comp1679minJ, comp2701minVal, comp2701minI, comp2701minJ);
    wire [11:0] comp2702minVal;
    wire [5:0] comp2702minI, comp2702minJ;
    Comparator comp2702(comp1680minVal, comp1680minI, comp1680minJ, comp1681minVal, comp1681minI, comp1681minJ, comp2702minVal, comp2702minI, comp2702minJ);
    wire [11:0] comp2703minVal;
    wire [5:0] comp2703minI, comp2703minJ;
    Comparator comp2703(comp1682minVal, comp1682minI, comp1682minJ, comp1683minVal, comp1683minI, comp1683minJ, comp2703minVal, comp2703minI, comp2703minJ);
    wire [11:0] comp2704minVal;
    wire [5:0] comp2704minI, comp2704minJ;
    Comparator comp2704(comp1684minVal, comp1684minI, comp1684minJ, comp1685minVal, comp1685minI, comp1685minJ, comp2704minVal, comp2704minI, comp2704minJ);
    wire [11:0] comp2705minVal;
    wire [5:0] comp2705minI, comp2705minJ;
    Comparator comp2705(comp1686minVal, comp1686minI, comp1686minJ, comp1687minVal, comp1687minI, comp1687minJ, comp2705minVal, comp2705minI, comp2705minJ);
    wire [11:0] comp2706minVal;
    wire [5:0] comp2706minI, comp2706minJ;
    Comparator comp2706(comp1688minVal, comp1688minI, comp1688minJ, comp1689minVal, comp1689minI, comp1689minJ, comp2706minVal, comp2706minI, comp2706minJ);
    wire [11:0] comp2707minVal;
    wire [5:0] comp2707minI, comp2707minJ;
    Comparator comp2707(comp1690minVal, comp1690minI, comp1690minJ, comp1691minVal, comp1691minI, comp1691minJ, comp2707minVal, comp2707minI, comp2707minJ);
    wire [11:0] comp2708minVal;
    wire [5:0] comp2708minI, comp2708minJ;
    Comparator comp2708(comp1692minVal, comp1692minI, comp1692minJ, comp1693minVal, comp1693minI, comp1693minJ, comp2708minVal, comp2708minI, comp2708minJ);
    wire [11:0] comp2709minVal;
    wire [5:0] comp2709minI, comp2709minJ;
    Comparator comp2709(comp1694minVal, comp1694minI, comp1694minJ, comp1695minVal, comp1695minI, comp1695minJ, comp2709minVal, comp2709minI, comp2709minJ);
    wire [11:0] comp2710minVal;
    wire [5:0] comp2710minI, comp2710minJ;
    Comparator comp2710(comp1696minVal, comp1696minI, comp1696minJ, comp1697minVal, comp1697minI, comp1697minJ, comp2710minVal, comp2710minI, comp2710minJ);
    wire [11:0] comp2711minVal;
    wire [5:0] comp2711minI, comp2711minJ;
    Comparator comp2711(comp1698minVal, comp1698minI, comp1698minJ, comp1699minVal, comp1699minI, comp1699minJ, comp2711minVal, comp2711minI, comp2711minJ);
    wire [11:0] comp2712minVal;
    wire [5:0] comp2712minI, comp2712minJ;
    Comparator comp2712(comp1700minVal, comp1700minI, comp1700minJ, comp1701minVal, comp1701minI, comp1701minJ, comp2712minVal, comp2712minI, comp2712minJ);
    wire [11:0] comp2713minVal;
    wire [5:0] comp2713minI, comp2713minJ;
    Comparator comp2713(comp1702minVal, comp1702minI, comp1702minJ, comp1703minVal, comp1703minI, comp1703minJ, comp2713minVal, comp2713minI, comp2713minJ);
    wire [11:0] comp2714minVal;
    wire [5:0] comp2714minI, comp2714minJ;
    Comparator comp2714(comp1704minVal, comp1704minI, comp1704minJ, comp1705minVal, comp1705minI, comp1705minJ, comp2714minVal, comp2714minI, comp2714minJ);
    wire [11:0] comp2715minVal;
    wire [5:0] comp2715minI, comp2715minJ;
    Comparator comp2715(comp1706minVal, comp1706minI, comp1706minJ, comp1707minVal, comp1707minI, comp1707minJ, comp2715minVal, comp2715minI, comp2715minJ);
    wire [11:0] comp2716minVal;
    wire [5:0] comp2716minI, comp2716minJ;
    Comparator comp2716(comp1708minVal, comp1708minI, comp1708minJ, comp1709minVal, comp1709minI, comp1709minJ, comp2716minVal, comp2716minI, comp2716minJ);
    wire [11:0] comp2717minVal;
    wire [5:0] comp2717minI, comp2717minJ;
    Comparator comp2717(comp1710minVal, comp1710minI, comp1710minJ, comp1711minVal, comp1711minI, comp1711minJ, comp2717minVal, comp2717minI, comp2717minJ);
    wire [11:0] comp2718minVal;
    wire [5:0] comp2718minI, comp2718minJ;
    Comparator comp2718(comp1712minVal, comp1712minI, comp1712minJ, comp1713minVal, comp1713minI, comp1713minJ, comp2718minVal, comp2718minI, comp2718minJ);
    wire [11:0] comp2719minVal;
    wire [5:0] comp2719minI, comp2719minJ;
    Comparator comp2719(comp1714minVal, comp1714minI, comp1714minJ, comp1715minVal, comp1715minI, comp1715minJ, comp2719minVal, comp2719minI, comp2719minJ);
    wire [11:0] comp2720minVal;
    wire [5:0] comp2720minI, comp2720minJ;
    Comparator comp2720(comp1716minVal, comp1716minI, comp1716minJ, comp1717minVal, comp1717minI, comp1717minJ, comp2720minVal, comp2720minI, comp2720minJ);
    wire [11:0] comp2721minVal;
    wire [5:0] comp2721minI, comp2721minJ;
    Comparator comp2721(comp1718minVal, comp1718minI, comp1718minJ, comp1719minVal, comp1719minI, comp1719minJ, comp2721minVal, comp2721minI, comp2721minJ);
    wire [11:0] comp2722minVal;
    wire [5:0] comp2722minI, comp2722minJ;
    Comparator comp2722(comp1720minVal, comp1720minI, comp1720minJ, comp1721minVal, comp1721minI, comp1721minJ, comp2722minVal, comp2722minI, comp2722minJ);
    wire [11:0] comp2723minVal;
    wire [5:0] comp2723minI, comp2723minJ;
    Comparator comp2723(comp1722minVal, comp1722minI, comp1722minJ, comp1723minVal, comp1723minI, comp1723minJ, comp2723minVal, comp2723minI, comp2723minJ);
    wire [11:0] comp2724minVal;
    wire [5:0] comp2724minI, comp2724minJ;
    Comparator comp2724(comp1724minVal, comp1724minI, comp1724minJ, comp1725minVal, comp1725minI, comp1725minJ, comp2724minVal, comp2724minI, comp2724minJ);
    wire [11:0] comp2725minVal;
    wire [5:0] comp2725minI, comp2725minJ;
    Comparator comp2725(comp1726minVal, comp1726minI, comp1726minJ, comp1727minVal, comp1727minI, comp1727minJ, comp2725minVal, comp2725minI, comp2725minJ);
    wire [11:0] comp2726minVal;
    wire [5:0] comp2726minI, comp2726minJ;
    Comparator comp2726(comp1728minVal, comp1728minI, comp1728minJ, comp1729minVal, comp1729minI, comp1729minJ, comp2726minVal, comp2726minI, comp2726minJ);
    wire [11:0] comp2727minVal;
    wire [5:0] comp2727minI, comp2727minJ;
    Comparator comp2727(comp1730minVal, comp1730minI, comp1730minJ, comp1731minVal, comp1731minI, comp1731minJ, comp2727minVal, comp2727minI, comp2727minJ);
    wire [11:0] comp2728minVal;
    wire [5:0] comp2728minI, comp2728minJ;
    Comparator comp2728(comp1732minVal, comp1732minI, comp1732minJ, comp1733minVal, comp1733minI, comp1733minJ, comp2728minVal, comp2728minI, comp2728minJ);
    wire [11:0] comp2729minVal;
    wire [5:0] comp2729minI, comp2729minJ;
    Comparator comp2729(comp1734minVal, comp1734minI, comp1734minJ, comp1735minVal, comp1735minI, comp1735minJ, comp2729minVal, comp2729minI, comp2729minJ);
    wire [11:0] comp2730minVal;
    wire [5:0] comp2730minI, comp2730minJ;
    Comparator comp2730(comp1736minVal, comp1736minI, comp1736minJ, comp1737minVal, comp1737minI, comp1737minJ, comp2730minVal, comp2730minI, comp2730minJ);
    wire [11:0] comp2731minVal;
    wire [5:0] comp2731minI, comp2731minJ;
    Comparator comp2731(comp1738minVal, comp1738minI, comp1738minJ, comp1739minVal, comp1739minI, comp1739minJ, comp2731minVal, comp2731minI, comp2731minJ);
    wire [11:0] comp2732minVal;
    wire [5:0] comp2732minI, comp2732minJ;
    Comparator comp2732(comp1740minVal, comp1740minI, comp1740minJ, comp1741minVal, comp1741minI, comp1741minJ, comp2732minVal, comp2732minI, comp2732minJ);
    wire [11:0] comp2733minVal;
    wire [5:0] comp2733minI, comp2733minJ;
    Comparator comp2733(comp1742minVal, comp1742minI, comp1742minJ, comp1743minVal, comp1743minI, comp1743minJ, comp2733minVal, comp2733minI, comp2733minJ);
    wire [11:0] comp2734minVal;
    wire [5:0] comp2734minI, comp2734minJ;
    Comparator comp2734(comp1744minVal, comp1744minI, comp1744minJ, comp1745minVal, comp1745minI, comp1745minJ, comp2734minVal, comp2734minI, comp2734minJ);
    wire [11:0] comp2735minVal;
    wire [5:0] comp2735minI, comp2735minJ;
    Comparator comp2735(comp1746minVal, comp1746minI, comp1746minJ, comp1747minVal, comp1747minI, comp1747minJ, comp2735minVal, comp2735minI, comp2735minJ);
    wire [11:0] comp2736minVal;
    wire [5:0] comp2736minI, comp2736minJ;
    Comparator comp2736(comp1748minVal, comp1748minI, comp1748minJ, comp1749minVal, comp1749minI, comp1749minJ, comp2736minVal, comp2736minI, comp2736minJ);
    wire [11:0] comp2737minVal;
    wire [5:0] comp2737minI, comp2737minJ;
    Comparator comp2737(comp1750minVal, comp1750minI, comp1750minJ, comp1751minVal, comp1751minI, comp1751minJ, comp2737minVal, comp2737minI, comp2737minJ);
    wire [11:0] comp2738minVal;
    wire [5:0] comp2738minI, comp2738minJ;
    Comparator comp2738(comp1752minVal, comp1752minI, comp1752minJ, comp1753minVal, comp1753minI, comp1753minJ, comp2738minVal, comp2738minI, comp2738minJ);
    wire [11:0] comp2739minVal;
    wire [5:0] comp2739minI, comp2739minJ;
    Comparator comp2739(comp1754minVal, comp1754minI, comp1754minJ, comp1755minVal, comp1755minI, comp1755minJ, comp2739minVal, comp2739minI, comp2739minJ);
    wire [11:0] comp2740minVal;
    wire [5:0] comp2740minI, comp2740minJ;
    Comparator comp2740(comp1756minVal, comp1756minI, comp1756minJ, comp1757minVal, comp1757minI, comp1757minJ, comp2740minVal, comp2740minI, comp2740minJ);
    wire [11:0] comp2741minVal;
    wire [5:0] comp2741minI, comp2741minJ;
    Comparator comp2741(comp1758minVal, comp1758minI, comp1758minJ, comp1759minVal, comp1759minI, comp1759minJ, comp2741minVal, comp2741minI, comp2741minJ);
    wire [11:0] comp2742minVal;
    wire [5:0] comp2742minI, comp2742minJ;
    Comparator comp2742(comp1760minVal, comp1760minI, comp1760minJ, comp1761minVal, comp1761minI, comp1761minJ, comp2742minVal, comp2742minI, comp2742minJ);
    wire [11:0] comp2743minVal;
    wire [5:0] comp2743minI, comp2743minJ;
    Comparator comp2743(comp1762minVal, comp1762minI, comp1762minJ, comp1763minVal, comp1763minI, comp1763minJ, comp2743minVal, comp2743minI, comp2743minJ);
    wire [11:0] comp2744minVal;
    wire [5:0] comp2744minI, comp2744minJ;
    Comparator comp2744(comp1764minVal, comp1764minI, comp1764minJ, comp1765minVal, comp1765minI, comp1765minJ, comp2744minVal, comp2744minI, comp2744minJ);
    wire [11:0] comp2745minVal;
    wire [5:0] comp2745minI, comp2745minJ;
    Comparator comp2745(comp1766minVal, comp1766minI, comp1766minJ, comp1767minVal, comp1767minI, comp1767minJ, comp2745minVal, comp2745minI, comp2745minJ);
    wire [11:0] comp2746minVal;
    wire [5:0] comp2746minI, comp2746minJ;
    Comparator comp2746(comp1768minVal, comp1768minI, comp1768minJ, comp1769minVal, comp1769minI, comp1769minJ, comp2746minVal, comp2746minI, comp2746minJ);
    wire [11:0] comp2747minVal;
    wire [5:0] comp2747minI, comp2747minJ;
    Comparator comp2747(comp1770minVal, comp1770minI, comp1770minJ, comp1771minVal, comp1771minI, comp1771minJ, comp2747minVal, comp2747minI, comp2747minJ);
    wire [11:0] comp2748minVal;
    wire [5:0] comp2748minI, comp2748minJ;
    Comparator comp2748(comp1772minVal, comp1772minI, comp1772minJ, comp1773minVal, comp1773minI, comp1773minJ, comp2748minVal, comp2748minI, comp2748minJ);
    wire [11:0] comp2749minVal;
    wire [5:0] comp2749minI, comp2749minJ;
    Comparator comp2749(comp1774minVal, comp1774minI, comp1774minJ, comp1775minVal, comp1775minI, comp1775minJ, comp2749minVal, comp2749minI, comp2749minJ);
    wire [11:0] comp2750minVal;
    wire [5:0] comp2750minI, comp2750minJ;
    Comparator comp2750(comp1776minVal, comp1776minI, comp1776minJ, comp1777minVal, comp1777minI, comp1777minJ, comp2750minVal, comp2750minI, comp2750minJ);
    wire [11:0] comp2751minVal;
    wire [5:0] comp2751minI, comp2751minJ;
    Comparator comp2751(comp1778minVal, comp1778minI, comp1778minJ, comp1779minVal, comp1779minI, comp1779minJ, comp2751minVal, comp2751minI, comp2751minJ);
    wire [11:0] comp2752minVal;
    wire [5:0] comp2752minI, comp2752minJ;
    Comparator comp2752(comp1780minVal, comp1780minI, comp1780minJ, comp1781minVal, comp1781minI, comp1781minJ, comp2752minVal, comp2752minI, comp2752minJ);
    wire [11:0] comp2753minVal;
    wire [5:0] comp2753minI, comp2753minJ;
    Comparator comp2753(comp1782minVal, comp1782minI, comp1782minJ, comp1783minVal, comp1783minI, comp1783minJ, comp2753minVal, comp2753minI, comp2753minJ);
    wire [11:0] comp2754minVal;
    wire [5:0] comp2754minI, comp2754minJ;
    Comparator comp2754(comp1784minVal, comp1784minI, comp1784minJ, comp1785minVal, comp1785minI, comp1785minJ, comp2754minVal, comp2754minI, comp2754minJ);
    wire [11:0] comp2755minVal;
    wire [5:0] comp2755minI, comp2755minJ;
    Comparator comp2755(comp1786minVal, comp1786minI, comp1786minJ, comp1787minVal, comp1787minI, comp1787minJ, comp2755minVal, comp2755minI, comp2755minJ);
    wire [11:0] comp2756minVal;
    wire [5:0] comp2756minI, comp2756minJ;
    Comparator comp2756(comp1788minVal, comp1788minI, comp1788minJ, comp1789minVal, comp1789minI, comp1789minJ, comp2756minVal, comp2756minI, comp2756minJ);
    wire [11:0] comp2757minVal;
    wire [5:0] comp2757minI, comp2757minJ;
    Comparator comp2757(comp1790minVal, comp1790minI, comp1790minJ, comp1791minVal, comp1791minI, comp1791minJ, comp2757minVal, comp2757minI, comp2757minJ);
    wire [11:0] comp2758minVal;
    wire [5:0] comp2758minI, comp2758minJ;
    Comparator comp2758(comp1792minVal, comp1792minI, comp1792minJ, comp1793minVal, comp1793minI, comp1793minJ, comp2758minVal, comp2758minI, comp2758minJ);
    wire [11:0] comp2759minVal;
    wire [5:0] comp2759minI, comp2759minJ;
    Comparator comp2759(comp1794minVal, comp1794minI, comp1794minJ, comp1795minVal, comp1795minI, comp1795minJ, comp2759minVal, comp2759minI, comp2759minJ);
    wire [11:0] comp2760minVal;
    wire [5:0] comp2760minI, comp2760minJ;
    Comparator comp2760(comp1796minVal, comp1796minI, comp1796minJ, comp1797minVal, comp1797minI, comp1797minJ, comp2760minVal, comp2760minI, comp2760minJ);
    wire [11:0] comp2761minVal;
    wire [5:0] comp2761minI, comp2761minJ;
    Comparator comp2761(comp1798minVal, comp1798minI, comp1798minJ, comp1799minVal, comp1799minI, comp1799minJ, comp2761minVal, comp2761minI, comp2761minJ);
    wire [11:0] comp2762minVal;
    wire [5:0] comp2762minI, comp2762minJ;
    Comparator comp2762(comp1800minVal, comp1800minI, comp1800minJ, comp1801minVal, comp1801minI, comp1801minJ, comp2762minVal, comp2762minI, comp2762minJ);
    wire [11:0] comp2763minVal;
    wire [5:0] comp2763minI, comp2763minJ;
    Comparator comp2763(comp1802minVal, comp1802minI, comp1802minJ, comp1803minVal, comp1803minI, comp1803minJ, comp2763minVal, comp2763minI, comp2763minJ);
    wire [11:0] comp2764minVal;
    wire [5:0] comp2764minI, comp2764minJ;
    Comparator comp2764(comp1804minVal, comp1804minI, comp1804minJ, comp1805minVal, comp1805minI, comp1805minJ, comp2764minVal, comp2764minI, comp2764minJ);
    wire [11:0] comp2765minVal;
    wire [5:0] comp2765minI, comp2765minJ;
    Comparator comp2765(comp1806minVal, comp1806minI, comp1806minJ, comp1807minVal, comp1807minI, comp1807minJ, comp2765minVal, comp2765minI, comp2765minJ);
    wire [11:0] comp2766minVal;
    wire [5:0] comp2766minI, comp2766minJ;
    Comparator comp2766(comp1808minVal, comp1808minI, comp1808minJ, comp1809minVal, comp1809minI, comp1809minJ, comp2766minVal, comp2766minI, comp2766minJ);
    wire [11:0] comp2767minVal;
    wire [5:0] comp2767minI, comp2767minJ;
    Comparator comp2767(comp1810minVal, comp1810minI, comp1810minJ, comp1811minVal, comp1811minI, comp1811minJ, comp2767minVal, comp2767minI, comp2767minJ);
    wire [11:0] comp2768minVal;
    wire [5:0] comp2768minI, comp2768minJ;
    Comparator comp2768(comp1812minVal, comp1812minI, comp1812minJ, comp1813minVal, comp1813minI, comp1813minJ, comp2768minVal, comp2768minI, comp2768minJ);
    wire [11:0] comp2769minVal;
    wire [5:0] comp2769minI, comp2769minJ;
    Comparator comp2769(comp1814minVal, comp1814minI, comp1814minJ, comp1815minVal, comp1815minI, comp1815minJ, comp2769minVal, comp2769minI, comp2769minJ);
    wire [11:0] comp2770minVal;
    wire [5:0] comp2770minI, comp2770minJ;
    Comparator comp2770(comp1816minVal, comp1816minI, comp1816minJ, comp1817minVal, comp1817minI, comp1817minJ, comp2770minVal, comp2770minI, comp2770minJ);
    wire [11:0] comp2771minVal;
    wire [5:0] comp2771minI, comp2771minJ;
    Comparator comp2771(comp1818minVal, comp1818minI, comp1818minJ, comp1819minVal, comp1819minI, comp1819minJ, comp2771minVal, comp2771minI, comp2771minJ);
    wire [11:0] comp2772minVal;
    wire [5:0] comp2772minI, comp2772minJ;
    Comparator comp2772(comp1820minVal, comp1820minI, comp1820minJ, comp1821minVal, comp1821minI, comp1821minJ, comp2772minVal, comp2772minI, comp2772minJ);
    wire [11:0] comp2773minVal;
    wire [5:0] comp2773minI, comp2773minJ;
    Comparator comp2773(comp1822minVal, comp1822minI, comp1822minJ, comp1823minVal, comp1823minI, comp1823minJ, comp2773minVal, comp2773minI, comp2773minJ);
    wire [11:0] comp2774minVal;
    wire [5:0] comp2774minI, comp2774minJ;
    Comparator comp2774(comp1824minVal, comp1824minI, comp1824minJ, comp1825minVal, comp1825minI, comp1825minJ, comp2774minVal, comp2774minI, comp2774minJ);
    wire [11:0] comp2775minVal;
    wire [5:0] comp2775minI, comp2775minJ;
    Comparator comp2775(comp1826minVal, comp1826minI, comp1826minJ, comp1827minVal, comp1827minI, comp1827minJ, comp2775minVal, comp2775minI, comp2775minJ);
    wire [11:0] comp2776minVal;
    wire [5:0] comp2776minI, comp2776minJ;
    Comparator comp2776(comp1828minVal, comp1828minI, comp1828minJ, comp1829minVal, comp1829minI, comp1829minJ, comp2776minVal, comp2776minI, comp2776minJ);
    wire [11:0] comp2777minVal;
    wire [5:0] comp2777minI, comp2777minJ;
    Comparator comp2777(comp1830minVal, comp1830minI, comp1830minJ, comp1831minVal, comp1831minI, comp1831minJ, comp2777minVal, comp2777minI, comp2777minJ);
    wire [11:0] comp2778minVal;
    wire [5:0] comp2778minI, comp2778minJ;
    Comparator comp2778(comp1832minVal, comp1832minI, comp1832minJ, comp1833minVal, comp1833minI, comp1833minJ, comp2778minVal, comp2778minI, comp2778minJ);
    wire [11:0] comp2779minVal;
    wire [5:0] comp2779minI, comp2779minJ;
    Comparator comp2779(comp1834minVal, comp1834minI, comp1834minJ, comp1835minVal, comp1835minI, comp1835minJ, comp2779minVal, comp2779minI, comp2779minJ);
    wire [11:0] comp2780minVal;
    wire [5:0] comp2780minI, comp2780minJ;
    Comparator comp2780(comp1836minVal, comp1836minI, comp1836minJ, comp1837minVal, comp1837minI, comp1837minJ, comp2780minVal, comp2780minI, comp2780minJ);
    wire [11:0] comp2781minVal;
    wire [5:0] comp2781minI, comp2781minJ;
    Comparator comp2781(comp1838minVal, comp1838minI, comp1838minJ, comp1839minVal, comp1839minI, comp1839minJ, comp2781minVal, comp2781minI, comp2781minJ);
    wire [11:0] comp2782minVal;
    wire [5:0] comp2782minI, comp2782minJ;
    Comparator comp2782(comp1840minVal, comp1840minI, comp1840minJ, comp1841minVal, comp1841minI, comp1841minJ, comp2782minVal, comp2782minI, comp2782minJ);
    wire [11:0] comp2783minVal;
    wire [5:0] comp2783minI, comp2783minJ;
    Comparator comp2783(comp1842minVal, comp1842minI, comp1842minJ, comp1843minVal, comp1843minI, comp1843minJ, comp2783minVal, comp2783minI, comp2783minJ);
    wire [11:0] comp2784minVal;
    wire [5:0] comp2784minI, comp2784minJ;
    Comparator comp2784(comp1844minVal, comp1844minI, comp1844minJ, comp1845minVal, comp1845minI, comp1845minJ, comp2784minVal, comp2784minI, comp2784minJ);
    wire [11:0] comp2785minVal;
    wire [5:0] comp2785minI, comp2785minJ;
    Comparator comp2785(comp1846minVal, comp1846minI, comp1846minJ, comp1847minVal, comp1847minI, comp1847minJ, comp2785minVal, comp2785minI, comp2785minJ);
    wire [11:0] comp2786minVal;
    wire [5:0] comp2786minI, comp2786minJ;
    Comparator comp2786(comp1848minVal, comp1848minI, comp1848minJ, comp1849minVal, comp1849minI, comp1849minJ, comp2786minVal, comp2786minI, comp2786minJ);
    wire [11:0] comp2787minVal;
    wire [5:0] comp2787minI, comp2787minJ;
    Comparator comp2787(comp1850minVal, comp1850minI, comp1850minJ, comp1851minVal, comp1851minI, comp1851minJ, comp2787minVal, comp2787minI, comp2787minJ);
    wire [11:0] comp2788minVal;
    wire [5:0] comp2788minI, comp2788minJ;
    Comparator comp2788(comp1852minVal, comp1852minI, comp1852minJ, comp1853minVal, comp1853minI, comp1853minJ, comp2788minVal, comp2788minI, comp2788minJ);
    wire [11:0] comp2789minVal;
    wire [5:0] comp2789minI, comp2789minJ;
    Comparator comp2789(comp1854minVal, comp1854minI, comp1854minJ, comp1855minVal, comp1855minI, comp1855minJ, comp2789minVal, comp2789minI, comp2789minJ);
    wire [11:0] comp2790minVal;
    wire [5:0] comp2790minI, comp2790minJ;
    Comparator comp2790(comp1856minVal, comp1856minI, comp1856minJ, comp1857minVal, comp1857minI, comp1857minJ, comp2790minVal, comp2790minI, comp2790minJ);
    wire [11:0] comp2791minVal;
    wire [5:0] comp2791minI, comp2791minJ;
    Comparator comp2791(comp1858minVal, comp1858minI, comp1858minJ, comp1859minVal, comp1859minI, comp1859minJ, comp2791minVal, comp2791minI, comp2791minJ);
    wire [11:0] comp2792minVal;
    wire [5:0] comp2792minI, comp2792minJ;
    Comparator comp2792(comp1860minVal, comp1860minI, comp1860minJ, comp1861minVal, comp1861minI, comp1861minJ, comp2792minVal, comp2792minI, comp2792minJ);
    wire [11:0] comp2793minVal;
    wire [5:0] comp2793minI, comp2793minJ;
    assign comp2793minVal = 4095;
    assign comp2793minI = 0;
    assign comp2793minJ = 0;
    wire [11:0] comp2794minVal;
    wire [5:0] comp2794minI, comp2794minJ;
    Comparator comp2794(comp1862minVal, comp1862minI, comp1862minJ, comp1863minVal, comp1863minI, comp1863minJ, comp2794minVal, comp2794minI, comp2794minJ);
    wire [11:0] comp2795minVal;
    wire [5:0] comp2795minI, comp2795minJ;
    Comparator comp2795(comp1864minVal, comp1864minI, comp1864minJ, comp1865minVal, comp1865minI, comp1865minJ, comp2795minVal, comp2795minI, comp2795minJ);
    wire [11:0] comp2796minVal;
    wire [5:0] comp2796minI, comp2796minJ;
    Comparator comp2796(comp1866minVal, comp1866minI, comp1866minJ, comp1867minVal, comp1867minI, comp1867minJ, comp2796minVal, comp2796minI, comp2796minJ);
    wire [11:0] comp2797minVal;
    wire [5:0] comp2797minI, comp2797minJ;
    Comparator comp2797(comp1868minVal, comp1868minI, comp1868minJ, comp1869minVal, comp1869minI, comp1869minJ, comp2797minVal, comp2797minI, comp2797minJ);
    wire [11:0] comp2798minVal;
    wire [5:0] comp2798minI, comp2798minJ;
    Comparator comp2798(comp1870minVal, comp1870minI, comp1870minJ, comp1871minVal, comp1871minI, comp1871minJ, comp2798minVal, comp2798minI, comp2798minJ);
    wire [11:0] comp2799minVal;
    wire [5:0] comp2799minI, comp2799minJ;
    Comparator comp2799(comp1872minVal, comp1872minI, comp1872minJ, comp1873minVal, comp1873minI, comp1873minJ, comp2799minVal, comp2799minI, comp2799minJ);
    wire [11:0] comp2800minVal;
    wire [5:0] comp2800minI, comp2800minJ;
    Comparator comp2800(comp1874minVal, comp1874minI, comp1874minJ, comp1875minVal, comp1875minI, comp1875minJ, comp2800minVal, comp2800minI, comp2800minJ);
    wire [11:0] comp2801minVal;
    wire [5:0] comp2801minI, comp2801minJ;
    Comparator comp2801(comp1876minVal, comp1876minI, comp1876minJ, comp1877minVal, comp1877minI, comp1877minJ, comp2801minVal, comp2801minI, comp2801minJ);
    wire [11:0] comp2802minVal;
    wire [5:0] comp2802minI, comp2802minJ;
    Comparator comp2802(comp1878minVal, comp1878minI, comp1878minJ, comp1879minVal, comp1879minI, comp1879minJ, comp2802minVal, comp2802minI, comp2802minJ);
    wire [11:0] comp2803minVal;
    wire [5:0] comp2803minI, comp2803minJ;
    Comparator comp2803(comp1880minVal, comp1880minI, comp1880minJ, comp1881minVal, comp1881minI, comp1881minJ, comp2803minVal, comp2803minI, comp2803minJ);
    wire [11:0] comp2804minVal;
    wire [5:0] comp2804minI, comp2804minJ;
    Comparator comp2804(comp1882minVal, comp1882minI, comp1882minJ, comp1883minVal, comp1883minI, comp1883minJ, comp2804minVal, comp2804minI, comp2804minJ);
    wire [11:0] comp2805minVal;
    wire [5:0] comp2805minI, comp2805minJ;
    Comparator comp2805(comp1884minVal, comp1884minI, comp1884minJ, comp1885minVal, comp1885minI, comp1885minJ, comp2805minVal, comp2805minI, comp2805minJ);
    wire [11:0] comp2806minVal;
    wire [5:0] comp2806minI, comp2806minJ;
    Comparator comp2806(comp1886minVal, comp1886minI, comp1886minJ, comp1887minVal, comp1887minI, comp1887minJ, comp2806minVal, comp2806minI, comp2806minJ);
    wire [11:0] comp2807minVal;
    wire [5:0] comp2807minI, comp2807minJ;
    Comparator comp2807(comp1888minVal, comp1888minI, comp1888minJ, comp1889minVal, comp1889minI, comp1889minJ, comp2807minVal, comp2807minI, comp2807minJ);
    wire [11:0] comp2808minVal;
    wire [5:0] comp2808minI, comp2808minJ;
    Comparator comp2808(comp1890minVal, comp1890minI, comp1890minJ, comp1891minVal, comp1891minI, comp1891minJ, comp2808minVal, comp2808minI, comp2808minJ);
    wire [11:0] comp2809minVal;
    wire [5:0] comp2809minI, comp2809minJ;
    Comparator comp2809(comp1892minVal, comp1892minI, comp1892minJ, comp1893minVal, comp1893minI, comp1893minJ, comp2809minVal, comp2809minI, comp2809minJ);
    wire [11:0] comp2810minVal;
    wire [5:0] comp2810minI, comp2810minJ;
    Comparator comp2810(comp1894minVal, comp1894minI, comp1894minJ, comp1895minVal, comp1895minI, comp1895minJ, comp2810minVal, comp2810minI, comp2810minJ);
    wire [11:0] comp2811minVal;
    wire [5:0] comp2811minI, comp2811minJ;
    Comparator comp2811(comp1896minVal, comp1896minI, comp1896minJ, comp1897minVal, comp1897minI, comp1897minJ, comp2811minVal, comp2811minI, comp2811minJ);
    wire [11:0] comp2812minVal;
    wire [5:0] comp2812minI, comp2812minJ;
    Comparator comp2812(comp1898minVal, comp1898minI, comp1898minJ, comp1899minVal, comp1899minI, comp1899minJ, comp2812minVal, comp2812minI, comp2812minJ);
    wire [11:0] comp2813minVal;
    wire [5:0] comp2813minI, comp2813minJ;
    Comparator comp2813(comp1900minVal, comp1900minI, comp1900minJ, comp1901minVal, comp1901minI, comp1901minJ, comp2813minVal, comp2813minI, comp2813minJ);
    wire [11:0] comp2814minVal;
    wire [5:0] comp2814minI, comp2814minJ;
    Comparator comp2814(comp1902minVal, comp1902minI, comp1902minJ, comp1903minVal, comp1903minI, comp1903minJ, comp2814minVal, comp2814minI, comp2814minJ);
    wire [11:0] comp2815minVal;
    wire [5:0] comp2815minI, comp2815minJ;
    Comparator comp2815(comp1904minVal, comp1904minI, comp1904minJ, comp1905minVal, comp1905minI, comp1905minJ, comp2815minVal, comp2815minI, comp2815minJ);
    wire [11:0] comp2816minVal;
    wire [5:0] comp2816minI, comp2816minJ;
    Comparator comp2816(comp1906minVal, comp1906minI, comp1906minJ, comp1907minVal, comp1907minI, comp1907minJ, comp2816minVal, comp2816minI, comp2816minJ);
    wire [11:0] comp2817minVal;
    wire [5:0] comp2817minI, comp2817minJ;
    Comparator comp2817(comp1908minVal, comp1908minI, comp1908minJ, comp1909minVal, comp1909minI, comp1909minJ, comp2817minVal, comp2817minI, comp2817minJ);
    wire [11:0] comp2818minVal;
    wire [5:0] comp2818minI, comp2818minJ;
    Comparator comp2818(comp1910minVal, comp1910minI, comp1910minJ, comp1911minVal, comp1911minI, comp1911minJ, comp2818minVal, comp2818minI, comp2818minJ);
    wire [11:0] comp2819minVal;
    wire [5:0] comp2819minI, comp2819minJ;
    Comparator comp2819(comp1912minVal, comp1912minI, comp1912minJ, comp1913minVal, comp1913minI, comp1913minJ, comp2819minVal, comp2819minI, comp2819minJ);
    wire [11:0] comp2820minVal;
    wire [5:0] comp2820minI, comp2820minJ;
    Comparator comp2820(comp1914minVal, comp1914minI, comp1914minJ, comp1915minVal, comp1915minI, comp1915minJ, comp2820minVal, comp2820minI, comp2820minJ);
    wire [11:0] comp2821minVal;
    wire [5:0] comp2821minI, comp2821minJ;
    Comparator comp2821(comp1916minVal, comp1916minI, comp1916minJ, comp1917minVal, comp1917minI, comp1917minJ, comp2821minVal, comp2821minI, comp2821minJ);
    wire [11:0] comp2822minVal;
    wire [5:0] comp2822minI, comp2822minJ;
    Comparator comp2822(comp1918minVal, comp1918minI, comp1918minJ, comp1919minVal, comp1919minI, comp1919minJ, comp2822minVal, comp2822minI, comp2822minJ);
    wire [11:0] comp2823minVal;
    wire [5:0] comp2823minI, comp2823minJ;
    Comparator comp2823(comp1920minVal, comp1920minI, comp1920minJ, comp1921minVal, comp1921minI, comp1921minJ, comp2823minVal, comp2823minI, comp2823minJ);
    wire [11:0] comp2824minVal;
    wire [5:0] comp2824minI, comp2824minJ;
    Comparator comp2824(comp1922minVal, comp1922minI, comp1922minJ, comp1923minVal, comp1923minI, comp1923minJ, comp2824minVal, comp2824minI, comp2824minJ);
    wire [11:0] comp2825minVal;
    wire [5:0] comp2825minI, comp2825minJ;
    Comparator comp2825(comp1924minVal, comp1924minI, comp1924minJ, comp1925minVal, comp1925minI, comp1925minJ, comp2825minVal, comp2825minI, comp2825minJ);
    wire [11:0] comp2826minVal;
    wire [5:0] comp2826minI, comp2826minJ;
    Comparator comp2826(comp1926minVal, comp1926minI, comp1926minJ, comp1927minVal, comp1927minI, comp1927minJ, comp2826minVal, comp2826minI, comp2826minJ);
    wire [11:0] comp2827minVal;
    wire [5:0] comp2827minI, comp2827minJ;
    Comparator comp2827(comp1928minVal, comp1928minI, comp1928minJ, comp1929minVal, comp1929minI, comp1929minJ, comp2827minVal, comp2827minI, comp2827minJ);
    wire [11:0] comp2828minVal;
    wire [5:0] comp2828minI, comp2828minJ;
    Comparator comp2828(comp1930minVal, comp1930minI, comp1930minJ, comp1931minVal, comp1931minI, comp1931minJ, comp2828minVal, comp2828minI, comp2828minJ);
    wire [11:0] comp2829minVal;
    wire [5:0] comp2829minI, comp2829minJ;
    Comparator comp2829(comp1932minVal, comp1932minI, comp1932minJ, comp1933minVal, comp1933minI, comp1933minJ, comp2829minVal, comp2829minI, comp2829minJ);
    wire [11:0] comp2830minVal;
    wire [5:0] comp2830minI, comp2830minJ;
    Comparator comp2830(comp1934minVal, comp1934minI, comp1934minJ, comp1935minVal, comp1935minI, comp1935minJ, comp2830minVal, comp2830minI, comp2830minJ);
    wire [11:0] comp2831minVal;
    wire [5:0] comp2831minI, comp2831minJ;
    Comparator comp2831(comp1936minVal, comp1936minI, comp1936minJ, comp1937minVal, comp1937minI, comp1937minJ, comp2831minVal, comp2831minI, comp2831minJ);
    wire [11:0] comp2832minVal;
    wire [5:0] comp2832minI, comp2832minJ;
    Comparator comp2832(comp1938minVal, comp1938minI, comp1938minJ, comp1939minVal, comp1939minI, comp1939minJ, comp2832minVal, comp2832minI, comp2832minJ);
    wire [11:0] comp2833minVal;
    wire [5:0] comp2833minI, comp2833minJ;
    Comparator comp2833(comp1940minVal, comp1940minI, comp1940minJ, comp1941minVal, comp1941minI, comp1941minJ, comp2833minVal, comp2833minI, comp2833minJ);
    wire [11:0] comp2834minVal;
    wire [5:0] comp2834minI, comp2834minJ;
    Comparator comp2834(comp1942minVal, comp1942minI, comp1942minJ, comp1943minVal, comp1943minI, comp1943minJ, comp2834minVal, comp2834minI, comp2834minJ);
    wire [11:0] comp2835minVal;
    wire [5:0] comp2835minI, comp2835minJ;
    Comparator comp2835(comp1944minVal, comp1944minI, comp1944minJ, comp1945minVal, comp1945minI, comp1945minJ, comp2835minVal, comp2835minI, comp2835minJ);
    wire [11:0] comp2836minVal;
    wire [5:0] comp2836minI, comp2836minJ;
    Comparator comp2836(comp1946minVal, comp1946minI, comp1946minJ, comp1947minVal, comp1947minI, comp1947minJ, comp2836minVal, comp2836minI, comp2836minJ);
    wire [11:0] comp2837minVal;
    wire [5:0] comp2837minI, comp2837minJ;
    Comparator comp2837(comp1948minVal, comp1948minI, comp1948minJ, comp1949minVal, comp1949minI, comp1949minJ, comp2837minVal, comp2837minI, comp2837minJ);
    wire [11:0] comp2838minVal;
    wire [5:0] comp2838minI, comp2838minJ;
    Comparator comp2838(comp1950minVal, comp1950minI, comp1950minJ, comp1951minVal, comp1951minI, comp1951minJ, comp2838minVal, comp2838minI, comp2838minJ);
    wire [11:0] comp2839minVal;
    wire [5:0] comp2839minI, comp2839minJ;
    Comparator comp2839(comp1952minVal, comp1952minI, comp1952minJ, comp1953minVal, comp1953minI, comp1953minJ, comp2839minVal, comp2839minI, comp2839minJ);
    wire [11:0] comp2840minVal;
    wire [5:0] comp2840minI, comp2840minJ;
    Comparator comp2840(comp1954minVal, comp1954minI, comp1954minJ, comp1955minVal, comp1955minI, comp1955minJ, comp2840minVal, comp2840minI, comp2840minJ);
    wire [11:0] comp2841minVal;
    wire [5:0] comp2841minI, comp2841minJ;
    Comparator comp2841(comp1956minVal, comp1956minI, comp1956minJ, comp1957minVal, comp1957minI, comp1957minJ, comp2841minVal, comp2841minI, comp2841minJ);
    wire [11:0] comp2842minVal;
    wire [5:0] comp2842minI, comp2842minJ;
    Comparator comp2842(comp1958minVal, comp1958minI, comp1958minJ, comp1959minVal, comp1959minI, comp1959minJ, comp2842minVal, comp2842minI, comp2842minJ);
    wire [11:0] comp2843minVal;
    wire [5:0] comp2843minI, comp2843minJ;
    Comparator comp2843(comp1960minVal, comp1960minI, comp1960minJ, comp1961minVal, comp1961minI, comp1961minJ, comp2843minVal, comp2843minI, comp2843minJ);
    wire [11:0] comp2844minVal;
    wire [5:0] comp2844minI, comp2844minJ;
    Comparator comp2844(comp1962minVal, comp1962minI, comp1962minJ, comp1963minVal, comp1963minI, comp1963minJ, comp2844minVal, comp2844minI, comp2844minJ);
    wire [11:0] comp2845minVal;
    wire [5:0] comp2845minI, comp2845minJ;
    Comparator comp2845(comp1964minVal, comp1964minI, comp1964minJ, comp1965minVal, comp1965minI, comp1965minJ, comp2845minVal, comp2845minI, comp2845minJ);
    wire [11:0] comp2846minVal;
    wire [5:0] comp2846minI, comp2846minJ;
    Comparator comp2846(comp1966minVal, comp1966minI, comp1966minJ, comp1967minVal, comp1967minI, comp1967minJ, comp2846minVal, comp2846minI, comp2846minJ);
    wire [11:0] comp2847minVal;
    wire [5:0] comp2847minI, comp2847minJ;
    Comparator comp2847(comp1968minVal, comp1968minI, comp1968minJ, comp1969minVal, comp1969minI, comp1969minJ, comp2847minVal, comp2847minI, comp2847minJ);
    wire [11:0] comp2848minVal;
    wire [5:0] comp2848minI, comp2848minJ;
    Comparator comp2848(comp1970minVal, comp1970minI, comp1970minJ, comp1971minVal, comp1971minI, comp1971minJ, comp2848minVal, comp2848minI, comp2848minJ);
    wire [11:0] comp2849minVal;
    wire [5:0] comp2849minI, comp2849minJ;
    Comparator comp2849(comp1972minVal, comp1972minI, comp1972minJ, comp1973minVal, comp1973minI, comp1973minJ, comp2849minVal, comp2849minI, comp2849minJ);
    wire [11:0] comp2850minVal;
    wire [5:0] comp2850minI, comp2850minJ;
    Comparator comp2850(comp1974minVal, comp1974minI, comp1974minJ, comp1975minVal, comp1975minI, comp1975minJ, comp2850minVal, comp2850minI, comp2850minJ);
    wire [11:0] comp2851minVal;
    wire [5:0] comp2851minI, comp2851minJ;
    Comparator comp2851(comp1976minVal, comp1976minI, comp1976minJ, comp1977minVal, comp1977minI, comp1977minJ, comp2851minVal, comp2851minI, comp2851minJ);
    wire [11:0] comp2852minVal;
    wire [5:0] comp2852minI, comp2852minJ;
    Comparator comp2852(comp1978minVal, comp1978minI, comp1978minJ, comp1979minVal, comp1979minI, comp1979minJ, comp2852minVal, comp2852minI, comp2852minJ);
    wire [11:0] comp2853minVal;
    wire [5:0] comp2853minI, comp2853minJ;
    Comparator comp2853(comp1980minVal, comp1980minI, comp1980minJ, comp1981minVal, comp1981minI, comp1981minJ, comp2853minVal, comp2853minI, comp2853minJ);
    wire [11:0] comp2854minVal;
    wire [5:0] comp2854minI, comp2854minJ;
    Comparator comp2854(comp1982minVal, comp1982minI, comp1982minJ, comp1983minVal, comp1983minI, comp1983minJ, comp2854minVal, comp2854minI, comp2854minJ);
    wire [11:0] comp2855minVal;
    wire [5:0] comp2855minI, comp2855minJ;
    Comparator comp2855(comp1984minVal, comp1984minI, comp1984minJ, comp1985minVal, comp1985minI, comp1985minJ, comp2855minVal, comp2855minI, comp2855minJ);
    wire [11:0] comp2856minVal;
    wire [5:0] comp2856minI, comp2856minJ;
    Comparator comp2856(comp1986minVal, comp1986minI, comp1986minJ, comp1987minVal, comp1987minI, comp1987minJ, comp2856minVal, comp2856minI, comp2856minJ);
    wire [11:0] comp2857minVal;
    wire [5:0] comp2857minI, comp2857minJ;
    Comparator comp2857(comp1988minVal, comp1988minI, comp1988minJ, comp1989minVal, comp1989minI, comp1989minJ, comp2857minVal, comp2857minI, comp2857minJ);
    wire [11:0] comp2858minVal;
    wire [5:0] comp2858minI, comp2858minJ;
    Comparator comp2858(comp1990minVal, comp1990minI, comp1990minJ, comp1991minVal, comp1991minI, comp1991minJ, comp2858minVal, comp2858minI, comp2858minJ);
    wire [11:0] comp2859minVal;
    wire [5:0] comp2859minI, comp2859minJ;
    Comparator comp2859(comp1992minVal, comp1992minI, comp1992minJ, comp1993minVal, comp1993minI, comp1993minJ, comp2859minVal, comp2859minI, comp2859minJ);
    wire [11:0] comp2860minVal;
    wire [5:0] comp2860minI, comp2860minJ;
    Comparator comp2860(comp1994minVal, comp1994minI, comp1994minJ, comp1995minVal, comp1995minI, comp1995minJ, comp2860minVal, comp2860minI, comp2860minJ);
    wire [11:0] comp2861minVal;
    wire [5:0] comp2861minI, comp2861minJ;
    Comparator comp2861(comp1996minVal, comp1996minI, comp1996minJ, comp1997minVal, comp1997minI, comp1997minJ, comp2861minVal, comp2861minI, comp2861minJ);
    wire [11:0] comp2862minVal;
    wire [5:0] comp2862minI, comp2862minJ;
    Comparator comp2862(comp1998minVal, comp1998minI, comp1998minJ, comp1999minVal, comp1999minI, comp1999minJ, comp2862minVal, comp2862minI, comp2862minJ);
    wire [11:0] comp2863minVal;
    wire [5:0] comp2863minI, comp2863minJ;
    Comparator comp2863(comp2000minVal, comp2000minI, comp2000minJ, comp2001minVal, comp2001minI, comp2001minJ, comp2863minVal, comp2863minI, comp2863minJ);
    wire [11:0] comp2864minVal;
    wire [5:0] comp2864minI, comp2864minJ;
    Comparator comp2864(comp2002minVal, comp2002minI, comp2002minJ, comp2003minVal, comp2003minI, comp2003minJ, comp2864minVal, comp2864minI, comp2864minJ);
    wire [11:0] comp2865minVal;
    wire [5:0] comp2865minI, comp2865minJ;
    Comparator comp2865(comp2004minVal, comp2004minI, comp2004minJ, comp2005minVal, comp2005minI, comp2005minJ, comp2865minVal, comp2865minI, comp2865minJ);
    wire [11:0] comp2866minVal;
    wire [5:0] comp2866minI, comp2866minJ;
    Comparator comp2866(comp2006minVal, comp2006minI, comp2006minJ, comp2007minVal, comp2007minI, comp2007minJ, comp2866minVal, comp2866minI, comp2866minJ);
    wire [11:0] comp2867minVal;
    wire [5:0] comp2867minI, comp2867minJ;
    Comparator comp2867(comp2008minVal, comp2008minI, comp2008minJ, comp2009minVal, comp2009minI, comp2009minJ, comp2867minVal, comp2867minI, comp2867minJ);
    wire [11:0] comp2868minVal;
    wire [5:0] comp2868minI, comp2868minJ;
    Comparator comp2868(comp2010minVal, comp2010minI, comp2010minJ, comp2011minVal, comp2011minI, comp2011minJ, comp2868minVal, comp2868minI, comp2868minJ);
    wire [11:0] comp2869minVal;
    wire [5:0] comp2869minI, comp2869minJ;
    Comparator comp2869(comp2012minVal, comp2012minI, comp2012minJ, comp2013minVal, comp2013minI, comp2013minJ, comp2869minVal, comp2869minI, comp2869minJ);
    wire [11:0] comp2870minVal;
    wire [5:0] comp2870minI, comp2870minJ;
    Comparator comp2870(comp2014minVal, comp2014minI, comp2014minJ, comp2015minVal, comp2015minI, comp2015minJ, comp2870minVal, comp2870minI, comp2870minJ);
    wire [11:0] comp2871minVal;
    wire [5:0] comp2871minI, comp2871minJ;
    Comparator comp2871(comp2016minVal, comp2016minI, comp2016minJ, comp2017minVal, comp2017minI, comp2017minJ, comp2871minVal, comp2871minI, comp2871minJ);
    wire [11:0] comp2872minVal;
    wire [5:0] comp2872minI, comp2872minJ;
    Comparator comp2872(comp2018minVal, comp2018minI, comp2018minJ, comp2019minVal, comp2019minI, comp2019minJ, comp2872minVal, comp2872minI, comp2872minJ);
    wire [11:0] comp2873minVal;
    wire [5:0] comp2873minI, comp2873minJ;
    Comparator comp2873(comp2020minVal, comp2020minI, comp2020minJ, comp2021minVal, comp2021minI, comp2021minJ, comp2873minVal, comp2873minI, comp2873minJ);
    wire [11:0] comp2874minVal;
    wire [5:0] comp2874minI, comp2874minJ;
    Comparator comp2874(comp2022minVal, comp2022minI, comp2022minJ, comp2023minVal, comp2023minI, comp2023minJ, comp2874minVal, comp2874minI, comp2874minJ);
    wire [11:0] comp2875minVal;
    wire [5:0] comp2875minI, comp2875minJ;
    Comparator comp2875(comp2024minVal, comp2024minI, comp2024minJ, comp2025minVal, comp2025minI, comp2025minJ, comp2875minVal, comp2875minI, comp2875minJ);
    wire [11:0] comp2876minVal;
    wire [5:0] comp2876minI, comp2876minJ;
    Comparator comp2876(comp2026minVal, comp2026minI, comp2026minJ, comp2027minVal, comp2027minI, comp2027minJ, comp2876minVal, comp2876minI, comp2876minJ);
    wire [11:0] comp2877minVal;
    wire [5:0] comp2877minI, comp2877minJ;
    Comparator comp2877(comp2028minVal, comp2028minI, comp2028minJ, comp2029minVal, comp2029minI, comp2029minJ, comp2877minVal, comp2877minI, comp2877minJ);
    wire [11:0] comp2878minVal;
    wire [5:0] comp2878minI, comp2878minJ;
    Comparator comp2878(comp2030minVal, comp2030minI, comp2030minJ, comp2031minVal, comp2031minI, comp2031minJ, comp2878minVal, comp2878minI, comp2878minJ);
    wire [11:0] comp2879minVal;
    wire [5:0] comp2879minI, comp2879minJ;
    Comparator comp2879(comp2032minVal, comp2032minI, comp2032minJ, comp2033minVal, comp2033minI, comp2033minJ, comp2879minVal, comp2879minI, comp2879minJ);
    wire [11:0] comp2880minVal;
    wire [5:0] comp2880minI, comp2880minJ;
    Comparator comp2880(comp2034minVal, comp2034minI, comp2034minJ, comp2035minVal, comp2035minI, comp2035minJ, comp2880minVal, comp2880minI, comp2880minJ);
    wire [11:0] comp2881minVal;
    wire [5:0] comp2881minI, comp2881minJ;
    Comparator comp2881(comp2036minVal, comp2036minI, comp2036minJ, comp2037minVal, comp2037minI, comp2037minJ, comp2881minVal, comp2881minI, comp2881minJ);
    wire [11:0] comp2882minVal;
    wire [5:0] comp2882minI, comp2882minJ;
    Comparator comp2882(comp2038minVal, comp2038minI, comp2038minJ, comp2039minVal, comp2039minI, comp2039minJ, comp2882minVal, comp2882minI, comp2882minJ);
    wire [11:0] comp2883minVal;
    wire [5:0] comp2883minI, comp2883minJ;
    Comparator comp2883(comp2040minVal, comp2040minI, comp2040minJ, comp2041minVal, comp2041minI, comp2041minJ, comp2883minVal, comp2883minI, comp2883minJ);
    wire [11:0] comp2884minVal;
    wire [5:0] comp2884minI, comp2884minJ;
    Comparator comp2884(comp2042minVal, comp2042minI, comp2042minJ, comp2043minVal, comp2043minI, comp2043minJ, comp2884minVal, comp2884minI, comp2884minJ);
    wire [11:0] comp2885minVal;
    wire [5:0] comp2885minI, comp2885minJ;
    Comparator comp2885(comp2044minVal, comp2044minI, comp2044minJ, comp2045minVal, comp2045minI, comp2045minJ, comp2885minVal, comp2885minI, comp2885minJ);
    wire [11:0] comp2886minVal;
    wire [5:0] comp2886minI, comp2886minJ;
    Comparator comp2886(comp2046minVal, comp2046minI, comp2046minJ, comp2047minVal, comp2047minI, comp2047minJ, comp2886minVal, comp2886minI, comp2886minJ);
    wire [11:0] comp2887minVal;
    wire [5:0] comp2887minI, comp2887minJ;
    Comparator comp2887(comp2048minVal, comp2048minI, comp2048minJ, comp2049minVal, comp2049minI, comp2049minJ, comp2887minVal, comp2887minI, comp2887minJ);
    wire [11:0] comp2888minVal;
    wire [5:0] comp2888minI, comp2888minJ;
    Comparator comp2888(comp2050minVal, comp2050minI, comp2050minJ, comp2051minVal, comp2051minI, comp2051minJ, comp2888minVal, comp2888minI, comp2888minJ);
    wire [11:0] comp2889minVal;
    wire [5:0] comp2889minI, comp2889minJ;
    Comparator comp2889(comp2052minVal, comp2052minI, comp2052minJ, comp2053minVal, comp2053minI, comp2053minJ, comp2889minVal, comp2889minI, comp2889minJ);
    wire [11:0] comp2890minVal;
    wire [5:0] comp2890minI, comp2890minJ;
    Comparator comp2890(comp2054minVal, comp2054minI, comp2054minJ, comp2055minVal, comp2055minI, comp2055minJ, comp2890minVal, comp2890minI, comp2890minJ);
    wire [11:0] comp2891minVal;
    wire [5:0] comp2891minI, comp2891minJ;
    Comparator comp2891(comp2056minVal, comp2056minI, comp2056minJ, comp2057minVal, comp2057minI, comp2057minJ, comp2891minVal, comp2891minI, comp2891minJ);
    wire [11:0] comp2892minVal;
    wire [5:0] comp2892minI, comp2892minJ;
    Comparator comp2892(comp2058minVal, comp2058minI, comp2058minJ, comp2059minVal, comp2059minI, comp2059minJ, comp2892minVal, comp2892minI, comp2892minJ);
    wire [11:0] comp2893minVal;
    wire [5:0] comp2893minI, comp2893minJ;
    Comparator comp2893(comp2060minVal, comp2060minI, comp2060minJ, comp2061minVal, comp2061minI, comp2061minJ, comp2893minVal, comp2893minI, comp2893minJ);
    wire [11:0] comp2894minVal;
    wire [5:0] comp2894minI, comp2894minJ;
    Comparator comp2894(comp2062minVal, comp2062minI, comp2062minJ, comp2063minVal, comp2063minI, comp2063minJ, comp2894minVal, comp2894minI, comp2894minJ);
    wire [11:0] comp2895minVal;
    wire [5:0] comp2895minI, comp2895minJ;
    Comparator comp2895(comp2064minVal, comp2064minI, comp2064minJ, comp2065minVal, comp2065minI, comp2065minJ, comp2895minVal, comp2895minI, comp2895minJ);
    wire [11:0] comp2896minVal;
    wire [5:0] comp2896minI, comp2896minJ;
    Comparator comp2896(comp2066minVal, comp2066minI, comp2066minJ, comp2067minVal, comp2067minI, comp2067minJ, comp2896minVal, comp2896minI, comp2896minJ);
    wire [11:0] comp2897minVal;
    wire [5:0] comp2897minI, comp2897minJ;
    Comparator comp2897(comp2068minVal, comp2068minI, comp2068minJ, comp2069minVal, comp2069minI, comp2069minJ, comp2897minVal, comp2897minI, comp2897minJ);
    wire [11:0] comp2898minVal;
    wire [5:0] comp2898minI, comp2898minJ;
    Comparator comp2898(comp2070minVal, comp2070minI, comp2070minJ, comp2071minVal, comp2071minI, comp2071minJ, comp2898minVal, comp2898minI, comp2898minJ);
    wire [11:0] comp2899minVal;
    wire [5:0] comp2899minI, comp2899minJ;
    Comparator comp2899(comp2072minVal, comp2072minI, comp2072minJ, comp2073minVal, comp2073minI, comp2073minJ, comp2899minVal, comp2899minI, comp2899minJ);
    wire [11:0] comp2900minVal;
    wire [5:0] comp2900minI, comp2900minJ;
    Comparator comp2900(comp2074minVal, comp2074minI, comp2074minJ, comp2075minVal, comp2075minI, comp2075minJ, comp2900minVal, comp2900minI, comp2900minJ);
    wire [11:0] comp2901minVal;
    wire [5:0] comp2901minI, comp2901minJ;
    Comparator comp2901(comp2076minVal, comp2076minI, comp2076minJ, comp2077minVal, comp2077minI, comp2077minJ, comp2901minVal, comp2901minI, comp2901minJ);
    wire [11:0] comp2902minVal;
    wire [5:0] comp2902minI, comp2902minJ;
    Comparator comp2902(comp2078minVal, comp2078minI, comp2078minJ, comp2079minVal, comp2079minI, comp2079minJ, comp2902minVal, comp2902minI, comp2902minJ);
    wire [11:0] comp2903minVal;
    wire [5:0] comp2903minI, comp2903minJ;
    Comparator comp2903(comp2080minVal, comp2080minI, comp2080minJ, comp2081minVal, comp2081minI, comp2081minJ, comp2903minVal, comp2903minI, comp2903minJ);
    wire [11:0] comp2904minVal;
    wire [5:0] comp2904minI, comp2904minJ;
    Comparator comp2904(comp2082minVal, comp2082minI, comp2082minJ, comp2083minVal, comp2083minI, comp2083minJ, comp2904minVal, comp2904minI, comp2904minJ);
    wire [11:0] comp2905minVal;
    wire [5:0] comp2905minI, comp2905minJ;
    Comparator comp2905(comp2084minVal, comp2084minI, comp2084minJ, comp2085minVal, comp2085minI, comp2085minJ, comp2905minVal, comp2905minI, comp2905minJ);
    wire [11:0] comp2906minVal;
    wire [5:0] comp2906minI, comp2906minJ;
    Comparator comp2906(comp2086minVal, comp2086minI, comp2086minJ, comp2087minVal, comp2087minI, comp2087minJ, comp2906minVal, comp2906minI, comp2906minJ);
    wire [11:0] comp2907minVal;
    wire [5:0] comp2907minI, comp2907minJ;
    Comparator comp2907(comp2088minVal, comp2088minI, comp2088minJ, comp2089minVal, comp2089minI, comp2089minJ, comp2907minVal, comp2907minI, comp2907minJ);
    wire [11:0] comp2908minVal;
    wire [5:0] comp2908minI, comp2908minJ;
    Comparator comp2908(comp2090minVal, comp2090minI, comp2090minJ, comp2091minVal, comp2091minI, comp2091minJ, comp2908minVal, comp2908minI, comp2908minJ);
    wire [11:0] comp2909minVal;
    wire [5:0] comp2909minI, comp2909minJ;
    Comparator comp2909(comp2092minVal, comp2092minI, comp2092minJ, comp2093minVal, comp2093minI, comp2093minJ, comp2909minVal, comp2909minI, comp2909minJ);
    wire [11:0] comp2910minVal;
    wire [5:0] comp2910minI, comp2910minJ;
    Comparator comp2910(comp2094minVal, comp2094minI, comp2094minJ, comp2095minVal, comp2095minI, comp2095minJ, comp2910minVal, comp2910minI, comp2910minJ);
    wire [11:0] comp2911minVal;
    wire [5:0] comp2911minI, comp2911minJ;
    Comparator comp2911(comp2096minVal, comp2096minI, comp2096minJ, comp2097minVal, comp2097minI, comp2097minJ, comp2911minVal, comp2911minI, comp2911minJ);
    wire [11:0] comp2912minVal;
    wire [5:0] comp2912minI, comp2912minJ;
    Comparator comp2912(comp2098minVal, comp2098minI, comp2098minJ, comp2099minVal, comp2099minI, comp2099minJ, comp2912minVal, comp2912minI, comp2912minJ);
    wire [11:0] comp2913minVal;
    wire [5:0] comp2913minI, comp2913minJ;
    Comparator comp2913(comp2100minVal, comp2100minI, comp2100minJ, comp2101minVal, comp2101minI, comp2101minJ, comp2913minVal, comp2913minI, comp2913minJ);
    wire [11:0] comp2914minVal;
    wire [5:0] comp2914minI, comp2914minJ;
    Comparator comp2914(comp2102minVal, comp2102minI, comp2102minJ, comp2103minVal, comp2103minI, comp2103minJ, comp2914minVal, comp2914minI, comp2914minJ);
    wire [11:0] comp2915minVal;
    wire [5:0] comp2915minI, comp2915minJ;
    Comparator comp2915(comp2104minVal, comp2104minI, comp2104minJ, comp2105minVal, comp2105minI, comp2105minJ, comp2915minVal, comp2915minI, comp2915minJ);
    wire [11:0] comp2916minVal;
    wire [5:0] comp2916minI, comp2916minJ;
    Comparator comp2916(comp2106minVal, comp2106minI, comp2106minJ, comp2107minVal, comp2107minI, comp2107minJ, comp2916minVal, comp2916minI, comp2916minJ);
    wire [11:0] comp2917minVal;
    wire [5:0] comp2917minI, comp2917minJ;
    Comparator comp2917(comp2108minVal, comp2108minI, comp2108minJ, comp2109minVal, comp2109minI, comp2109minJ, comp2917minVal, comp2917minI, comp2917minJ);
    wire [11:0] comp2918minVal;
    wire [5:0] comp2918minI, comp2918minJ;
    Comparator comp2918(comp2110minVal, comp2110minI, comp2110minJ, comp2111minVal, comp2111minI, comp2111minJ, comp2918minVal, comp2918minI, comp2918minJ);
    wire [11:0] comp2919minVal;
    wire [5:0] comp2919minI, comp2919minJ;
    Comparator comp2919(comp2112minVal, comp2112minI, comp2112minJ, comp2113minVal, comp2113minI, comp2113minJ, comp2919minVal, comp2919minI, comp2919minJ);
    wire [11:0] comp2920minVal;
    wire [5:0] comp2920minI, comp2920minJ;
    Comparator comp2920(comp2114minVal, comp2114minI, comp2114minJ, comp2115minVal, comp2115minI, comp2115minJ, comp2920minVal, comp2920minI, comp2920minJ);
    wire [11:0] comp2921minVal;
    wire [5:0] comp2921minI, comp2921minJ;
    Comparator comp2921(comp2116minVal, comp2116minI, comp2116minJ, comp2117minVal, comp2117minI, comp2117minJ, comp2921minVal, comp2921minI, comp2921minJ);
    wire [11:0] comp2922minVal;
    wire [5:0] comp2922minI, comp2922minJ;
    Comparator comp2922(comp2118minVal, comp2118minI, comp2118minJ, comp2119minVal, comp2119minI, comp2119minJ, comp2922minVal, comp2922minI, comp2922minJ);
    wire [11:0] comp2923minVal;
    wire [5:0] comp2923minI, comp2923minJ;
    Comparator comp2923(comp2120minVal, comp2120minI, comp2120minJ, comp2121minVal, comp2121minI, comp2121minJ, comp2923minVal, comp2923minI, comp2923minJ);
    wire [11:0] comp2924minVal;
    wire [5:0] comp2924minI, comp2924minJ;
    Comparator comp2924(comp2122minVal, comp2122minI, comp2122minJ, comp2123minVal, comp2123minI, comp2123minJ, comp2924minVal, comp2924minI, comp2924minJ);
    wire [11:0] comp2925minVal;
    wire [5:0] comp2925minI, comp2925minJ;
    Comparator comp2925(comp2124minVal, comp2124minI, comp2124minJ, comp2125minVal, comp2125minI, comp2125minJ, comp2925minVal, comp2925minI, comp2925minJ);
    wire [11:0] comp2926minVal;
    wire [5:0] comp2926minI, comp2926minJ;
    Comparator comp2926(comp2126minVal, comp2126minI, comp2126minJ, comp2127minVal, comp2127minI, comp2127minJ, comp2926minVal, comp2926minI, comp2926minJ);
    wire [11:0] comp2927minVal;
    wire [5:0] comp2927minI, comp2927minJ;
    Comparator comp2927(comp2128minVal, comp2128minI, comp2128minJ, comp2129minVal, comp2129minI, comp2129minJ, comp2927minVal, comp2927minI, comp2927minJ);
    wire [11:0] comp2928minVal;
    wire [5:0] comp2928minI, comp2928minJ;
    Comparator comp2928(comp2130minVal, comp2130minI, comp2130minJ, comp2131minVal, comp2131minI, comp2131minJ, comp2928minVal, comp2928minI, comp2928minJ);
    wire [11:0] comp2929minVal;
    wire [5:0] comp2929minI, comp2929minJ;
    Comparator comp2929(comp2132minVal, comp2132minI, comp2132minJ, comp2133minVal, comp2133minI, comp2133minJ, comp2929minVal, comp2929minI, comp2929minJ);
    wire [11:0] comp2930minVal;
    wire [5:0] comp2930minI, comp2930minJ;
    Comparator comp2930(comp2134minVal, comp2134minI, comp2134minJ, comp2135minVal, comp2135minI, comp2135minJ, comp2930minVal, comp2930minI, comp2930minJ);
    wire [11:0] comp2931minVal;
    wire [5:0] comp2931minI, comp2931minJ;
    Comparator comp2931(comp2136minVal, comp2136minI, comp2136minJ, comp2137minVal, comp2137minI, comp2137minJ, comp2931minVal, comp2931minI, comp2931minJ);
    wire [11:0] comp2932minVal;
    wire [5:0] comp2932minI, comp2932minJ;
    Comparator comp2932(comp2138minVal, comp2138minI, comp2138minJ, comp2139minVal, comp2139minI, comp2139minJ, comp2932minVal, comp2932minI, comp2932minJ);
    wire [11:0] comp2933minVal;
    wire [5:0] comp2933minI, comp2933minJ;
    Comparator comp2933(comp2140minVal, comp2140minI, comp2140minJ, comp2141minVal, comp2141minI, comp2141minJ, comp2933minVal, comp2933minI, comp2933minJ);
    wire [11:0] comp2934minVal;
    wire [5:0] comp2934minI, comp2934minJ;
    Comparator comp2934(comp2142minVal, comp2142minI, comp2142minJ, comp2143minVal, comp2143minI, comp2143minJ, comp2934minVal, comp2934minI, comp2934minJ);
    wire [11:0] comp2935minVal;
    wire [5:0] comp2935minI, comp2935minJ;
    Comparator comp2935(comp2144minVal, comp2144minI, comp2144minJ, comp2145minVal, comp2145minI, comp2145minJ, comp2935minVal, comp2935minI, comp2935minJ);
    wire [11:0] comp2936minVal;
    wire [5:0] comp2936minI, comp2936minJ;
    Comparator comp2936(comp2146minVal, comp2146minI, comp2146minJ, comp2147minVal, comp2147minI, comp2147minJ, comp2936minVal, comp2936minI, comp2936minJ);
    wire [11:0] comp2937minVal;
    wire [5:0] comp2937minI, comp2937minJ;
    Comparator comp2937(comp2148minVal, comp2148minI, comp2148minJ, comp2149minVal, comp2149minI, comp2149minJ, comp2937minVal, comp2937minI, comp2937minJ);
    wire [11:0] comp2938minVal;
    wire [5:0] comp2938minI, comp2938minJ;
    Comparator comp2938(comp2150minVal, comp2150minI, comp2150minJ, comp2151minVal, comp2151minI, comp2151minJ, comp2938minVal, comp2938minI, comp2938minJ);
    wire [11:0] comp2939minVal;
    wire [5:0] comp2939minI, comp2939minJ;
    Comparator comp2939(comp2152minVal, comp2152minI, comp2152minJ, comp2153minVal, comp2153minI, comp2153minJ, comp2939minVal, comp2939minI, comp2939minJ);
    wire [11:0] comp2940minVal;
    wire [5:0] comp2940minI, comp2940minJ;
    Comparator comp2940(comp2154minVal, comp2154minI, comp2154minJ, comp2155minVal, comp2155minI, comp2155minJ, comp2940minVal, comp2940minI, comp2940minJ);
    wire [11:0] comp2941minVal;
    wire [5:0] comp2941minI, comp2941minJ;
    Comparator comp2941(comp2156minVal, comp2156minI, comp2156minJ, comp2157minVal, comp2157minI, comp2157minJ, comp2941minVal, comp2941minI, comp2941minJ);
    wire [11:0] comp2942minVal;
    wire [5:0] comp2942minI, comp2942minJ;
    Comparator comp2942(comp2158minVal, comp2158minI, comp2158minJ, comp2159minVal, comp2159minI, comp2159minJ, comp2942minVal, comp2942minI, comp2942minJ);
    wire [11:0] comp2943minVal;
    wire [5:0] comp2943minI, comp2943minJ;
    Comparator comp2943(comp2160minVal, comp2160minI, comp2160minJ, comp2161minVal, comp2161minI, comp2161minJ, comp2943minVal, comp2943minI, comp2943minJ);
    wire [11:0] comp2944minVal;
    wire [5:0] comp2944minI, comp2944minJ;
    Comparator comp2944(comp2162minVal, comp2162minI, comp2162minJ, comp2163minVal, comp2163minI, comp2163minJ, comp2944minVal, comp2944minI, comp2944minJ);
    wire [11:0] comp2945minVal;
    wire [5:0] comp2945minI, comp2945minJ;
    Comparator comp2945(comp2164minVal, comp2164minI, comp2164minJ, comp2165minVal, comp2165minI, comp2165minJ, comp2945minVal, comp2945minI, comp2945minJ);
    wire [11:0] comp2946minVal;
    wire [5:0] comp2946minI, comp2946minJ;
    Comparator comp2946(comp2166minVal, comp2166minI, comp2166minJ, comp2167minVal, comp2167minI, comp2167minJ, comp2946minVal, comp2946minI, comp2946minJ);
    wire [11:0] comp2947minVal;
    wire [5:0] comp2947minI, comp2947minJ;
    Comparator comp2947(comp2168minVal, comp2168minI, comp2168minJ, comp2169minVal, comp2169minI, comp2169minJ, comp2947minVal, comp2947minI, comp2947minJ);
    wire [11:0] comp2948minVal;
    wire [5:0] comp2948minI, comp2948minJ;
    Comparator comp2948(comp2170minVal, comp2170minI, comp2170minJ, comp2171minVal, comp2171minI, comp2171minJ, comp2948minVal, comp2948minI, comp2948minJ);
    wire [11:0] comp2949minVal;
    wire [5:0] comp2949minI, comp2949minJ;
    Comparator comp2949(comp2172minVal, comp2172minI, comp2172minJ, comp2173minVal, comp2173minI, comp2173minJ, comp2949minVal, comp2949minI, comp2949minJ);
    wire [11:0] comp2950minVal;
    wire [5:0] comp2950minI, comp2950minJ;
    Comparator comp2950(comp2174minVal, comp2174minI, comp2174minJ, comp2175minVal, comp2175minI, comp2175minJ, comp2950minVal, comp2950minI, comp2950minJ);
    wire [11:0] comp2951minVal;
    wire [5:0] comp2951minI, comp2951minJ;
    Comparator comp2951(comp2176minVal, comp2176minI, comp2176minJ, comp2177minVal, comp2177minI, comp2177minJ, comp2951minVal, comp2951minI, comp2951minJ);
    wire [11:0] comp2952minVal;
    wire [5:0] comp2952minI, comp2952minJ;
    Comparator comp2952(comp2178minVal, comp2178minI, comp2178minJ, comp2179minVal, comp2179minI, comp2179minJ, comp2952minVal, comp2952minI, comp2952minJ);
    wire [11:0] comp2953minVal;
    wire [5:0] comp2953minI, comp2953minJ;
    Comparator comp2953(comp2180minVal, comp2180minI, comp2180minJ, comp2181minVal, comp2181minI, comp2181minJ, comp2953minVal, comp2953minI, comp2953minJ);
    wire [11:0] comp2954minVal;
    wire [5:0] comp2954minI, comp2954minJ;
    Comparator comp2954(comp2182minVal, comp2182minI, comp2182minJ, comp2183minVal, comp2183minI, comp2183minJ, comp2954minVal, comp2954minI, comp2954minJ);
    wire [11:0] comp2955minVal;
    wire [5:0] comp2955minI, comp2955minJ;
    Comparator comp2955(comp2184minVal, comp2184minI, comp2184minJ, comp2185minVal, comp2185minI, comp2185minJ, comp2955minVal, comp2955minI, comp2955minJ);
    wire [11:0] comp2956minVal;
    wire [5:0] comp2956minI, comp2956minJ;
    Comparator comp2956(comp2186minVal, comp2186minI, comp2186minJ, comp2187minVal, comp2187minI, comp2187minJ, comp2956minVal, comp2956minI, comp2956minJ);
    wire [11:0] comp2957minVal;
    wire [5:0] comp2957minI, comp2957minJ;
    Comparator comp2957(comp2188minVal, comp2188minI, comp2188minJ, comp2189minVal, comp2189minI, comp2189minJ, comp2957minVal, comp2957minI, comp2957minJ);
    wire [11:0] comp2958minVal;
    wire [5:0] comp2958minI, comp2958minJ;
    Comparator comp2958(comp2190minVal, comp2190minI, comp2190minJ, comp2191minVal, comp2191minI, comp2191minJ, comp2958minVal, comp2958minI, comp2958minJ);
    wire [11:0] comp2959minVal;
    wire [5:0] comp2959minI, comp2959minJ;
    Comparator comp2959(comp2192minVal, comp2192minI, comp2192minJ, comp2193minVal, comp2193minI, comp2193minJ, comp2959minVal, comp2959minI, comp2959minJ);
    wire [11:0] comp2960minVal;
    wire [5:0] comp2960minI, comp2960minJ;
    Comparator comp2960(comp2194minVal, comp2194minI, comp2194minJ, comp2195minVal, comp2195minI, comp2195minJ, comp2960minVal, comp2960minI, comp2960minJ);
    wire [11:0] comp2961minVal;
    wire [5:0] comp2961minI, comp2961minJ;
    Comparator comp2961(comp2196minVal, comp2196minI, comp2196minJ, comp2197minVal, comp2197minI, comp2197minJ, comp2961minVal, comp2961minI, comp2961minJ);
    wire [11:0] comp2962minVal;
    wire [5:0] comp2962minI, comp2962minJ;
    Comparator comp2962(comp2198minVal, comp2198minI, comp2198minJ, comp2199minVal, comp2199minI, comp2199minJ, comp2962minVal, comp2962minI, comp2962minJ);
    wire [11:0] comp2963minVal;
    wire [5:0] comp2963minI, comp2963minJ;
    Comparator comp2963(comp2200minVal, comp2200minI, comp2200minJ, comp2201minVal, comp2201minI, comp2201minJ, comp2963minVal, comp2963minI, comp2963minJ);
    wire [11:0] comp2964minVal;
    wire [5:0] comp2964minI, comp2964minJ;
    Comparator comp2964(comp2202minVal, comp2202minI, comp2202minJ, comp2203minVal, comp2203minI, comp2203minJ, comp2964minVal, comp2964minI, comp2964minJ);
    wire [11:0] comp2965minVal;
    wire [5:0] comp2965minI, comp2965minJ;
    Comparator comp2965(comp2204minVal, comp2204minI, comp2204minJ, comp2205minVal, comp2205minI, comp2205minJ, comp2965minVal, comp2965minI, comp2965minJ);
    wire [11:0] comp2966minVal;
    wire [5:0] comp2966minI, comp2966minJ;
    Comparator comp2966(comp2206minVal, comp2206minI, comp2206minJ, comp2207minVal, comp2207minI, comp2207minJ, comp2966minVal, comp2966minI, comp2966minJ);
    wire [11:0] comp2967minVal;
    wire [5:0] comp2967minI, comp2967minJ;
    Comparator comp2967(comp2208minVal, comp2208minI, comp2208minJ, comp2209minVal, comp2209minI, comp2209minJ, comp2967minVal, comp2967minI, comp2967minJ);
    wire [11:0] comp2968minVal;
    wire [5:0] comp2968minI, comp2968minJ;
    Comparator comp2968(comp2210minVal, comp2210minI, comp2210minJ, comp2211minVal, comp2211minI, comp2211minJ, comp2968minVal, comp2968minI, comp2968minJ);
    wire [11:0] comp2969minVal;
    wire [5:0] comp2969minI, comp2969minJ;
    Comparator comp2969(comp2212minVal, comp2212minI, comp2212minJ, comp2213minVal, comp2213minI, comp2213minJ, comp2969minVal, comp2969minI, comp2969minJ);
    wire [11:0] comp2970minVal;
    wire [5:0] comp2970minI, comp2970minJ;
    Comparator comp2970(comp2214minVal, comp2214minI, comp2214minJ, comp2215minVal, comp2215minI, comp2215minJ, comp2970minVal, comp2970minI, comp2970minJ);
    wire [11:0] comp2971minVal;
    wire [5:0] comp2971minI, comp2971minJ;
    Comparator comp2971(comp2216minVal, comp2216minI, comp2216minJ, comp2217minVal, comp2217minI, comp2217minJ, comp2971minVal, comp2971minI, comp2971minJ);
    wire [11:0] comp2972minVal;
    wire [5:0] comp2972minI, comp2972minJ;
    Comparator comp2972(comp2218minVal, comp2218minI, comp2218minJ, comp2219minVal, comp2219minI, comp2219minJ, comp2972minVal, comp2972minI, comp2972minJ);
    wire [11:0] comp2973minVal;
    wire [5:0] comp2973minI, comp2973minJ;
    Comparator comp2973(comp2220minVal, comp2220minI, comp2220minJ, comp2221minVal, comp2221minI, comp2221minJ, comp2973minVal, comp2973minI, comp2973minJ);
    wire [11:0] comp2974minVal;
    wire [5:0] comp2974minI, comp2974minJ;
    Comparator comp2974(comp2222minVal, comp2222minI, comp2222minJ, comp2223minVal, comp2223minI, comp2223minJ, comp2974minVal, comp2974minI, comp2974minJ);
    wire [11:0] comp2975minVal;
    wire [5:0] comp2975minI, comp2975minJ;
    Comparator comp2975(comp2224minVal, comp2224minI, comp2224minJ, comp2225minVal, comp2225minI, comp2225minJ, comp2975minVal, comp2975minI, comp2975minJ);
    wire [11:0] comp2976minVal;
    wire [5:0] comp2976minI, comp2976minJ;
    Comparator comp2976(comp2226minVal, comp2226minI, comp2226minJ, comp2227minVal, comp2227minI, comp2227minJ, comp2976minVal, comp2976minI, comp2976minJ);
    wire [11:0] comp2977minVal;
    wire [5:0] comp2977minI, comp2977minJ;
    Comparator comp2977(comp2228minVal, comp2228minI, comp2228minJ, comp2229minVal, comp2229minI, comp2229minJ, comp2977minVal, comp2977minI, comp2977minJ);
    wire [11:0] comp2978minVal;
    wire [5:0] comp2978minI, comp2978minJ;
    Comparator comp2978(comp2230minVal, comp2230minI, comp2230minJ, comp2231minVal, comp2231minI, comp2231minJ, comp2978minVal, comp2978minI, comp2978minJ);
    wire [11:0] comp2979minVal;
    wire [5:0] comp2979minI, comp2979minJ;
    Comparator comp2979(comp2232minVal, comp2232minI, comp2232minJ, comp2233minVal, comp2233minI, comp2233minJ, comp2979minVal, comp2979minI, comp2979minJ);
    wire [11:0] comp2980minVal;
    wire [5:0] comp2980minI, comp2980minJ;
    Comparator comp2980(comp2234minVal, comp2234minI, comp2234minJ, comp2235minVal, comp2235minI, comp2235minJ, comp2980minVal, comp2980minI, comp2980minJ);
    wire [11:0] comp2981minVal;
    wire [5:0] comp2981minI, comp2981minJ;
    Comparator comp2981(comp2236minVal, comp2236minI, comp2236minJ, comp2237minVal, comp2237minI, comp2237minJ, comp2981minVal, comp2981minI, comp2981minJ);
    wire [11:0] comp2982minVal;
    wire [5:0] comp2982minI, comp2982minJ;
    Comparator comp2982(comp2238minVal, comp2238minI, comp2238minJ, comp2239minVal, comp2239minI, comp2239minJ, comp2982minVal, comp2982minI, comp2982minJ);
    wire [11:0] comp2983minVal;
    wire [5:0] comp2983minI, comp2983minJ;
    Comparator comp2983(comp2240minVal, comp2240minI, comp2240minJ, comp2241minVal, comp2241minI, comp2241minJ, comp2983minVal, comp2983minI, comp2983minJ);
    wire [11:0] comp2984minVal;
    wire [5:0] comp2984minI, comp2984minJ;
    Comparator comp2984(comp2242minVal, comp2242minI, comp2242minJ, comp2243minVal, comp2243minI, comp2243minJ, comp2984minVal, comp2984minI, comp2984minJ);
    wire [11:0] comp2985minVal;
    wire [5:0] comp2985minI, comp2985minJ;
    Comparator comp2985(comp2244minVal, comp2244minI, comp2244minJ, comp2245minVal, comp2245minI, comp2245minJ, comp2985minVal, comp2985minI, comp2985minJ);
    wire [11:0] comp2986minVal;
    wire [5:0] comp2986minI, comp2986minJ;
    Comparator comp2986(comp2246minVal, comp2246minI, comp2246minJ, comp2247minVal, comp2247minI, comp2247minJ, comp2986minVal, comp2986minI, comp2986minJ);
    wire [11:0] comp2987minVal;
    wire [5:0] comp2987minI, comp2987minJ;
    Comparator comp2987(comp2248minVal, comp2248minI, comp2248minJ, comp2249minVal, comp2249minI, comp2249minJ, comp2987minVal, comp2987minI, comp2987minJ);
    wire [11:0] comp2988minVal;
    wire [5:0] comp2988minI, comp2988minJ;
    Comparator comp2988(comp2250minVal, comp2250minI, comp2250minJ, comp2251minVal, comp2251minI, comp2251minJ, comp2988minVal, comp2988minI, comp2988minJ);
    wire [11:0] comp2989minVal;
    wire [5:0] comp2989minI, comp2989minJ;
    Comparator comp2989(comp2252minVal, comp2252minI, comp2252minJ, comp2253minVal, comp2253minI, comp2253minJ, comp2989minVal, comp2989minI, comp2989minJ);
    wire [11:0] comp2990minVal;
    wire [5:0] comp2990minI, comp2990minJ;
    Comparator comp2990(comp2254minVal, comp2254minI, comp2254minJ, comp2255minVal, comp2255minI, comp2255minJ, comp2990minVal, comp2990minI, comp2990minJ);
    wire [11:0] comp2991minVal;
    wire [5:0] comp2991minI, comp2991minJ;
    Comparator comp2991(comp2256minVal, comp2256minI, comp2256minJ, comp2257minVal, comp2257minI, comp2257minJ, comp2991minVal, comp2991minI, comp2991minJ);
    wire [11:0] comp2992minVal;
    wire [5:0] comp2992minI, comp2992minJ;
    Comparator comp2992(comp2258minVal, comp2258minI, comp2258minJ, comp2259minVal, comp2259minI, comp2259minJ, comp2992minVal, comp2992minI, comp2992minJ);
    wire [11:0] comp2993minVal;
    wire [5:0] comp2993minI, comp2993minJ;
    Comparator comp2993(comp2260minVal, comp2260minI, comp2260minJ, comp2261minVal, comp2261minI, comp2261minJ, comp2993minVal, comp2993minI, comp2993minJ);
    wire [11:0] comp2994minVal;
    wire [5:0] comp2994minI, comp2994minJ;
    Comparator comp2994(comp2262minVal, comp2262minI, comp2262minJ, comp2263minVal, comp2263minI, comp2263minJ, comp2994minVal, comp2994minI, comp2994minJ);
    wire [11:0] comp2995minVal;
    wire [5:0] comp2995minI, comp2995minJ;
    Comparator comp2995(comp2264minVal, comp2264minI, comp2264minJ, comp2265minVal, comp2265minI, comp2265minJ, comp2995minVal, comp2995minI, comp2995minJ);
    wire [11:0] comp2996minVal;
    wire [5:0] comp2996minI, comp2996minJ;
    Comparator comp2996(comp2266minVal, comp2266minI, comp2266minJ, comp2267minVal, comp2267minI, comp2267minJ, comp2996minVal, comp2996minI, comp2996minJ);
    wire [11:0] comp2997minVal;
    wire [5:0] comp2997minI, comp2997minJ;
    Comparator comp2997(comp2268minVal, comp2268minI, comp2268minJ, comp2269minVal, comp2269minI, comp2269minJ, comp2997minVal, comp2997minI, comp2997minJ);
    wire [11:0] comp2998minVal;
    wire [5:0] comp2998minI, comp2998minJ;
    Comparator comp2998(comp2270minVal, comp2270minI, comp2270minJ, comp2271minVal, comp2271minI, comp2271minJ, comp2998minVal, comp2998minI, comp2998minJ);
    wire [11:0] comp2999minVal;
    wire [5:0] comp2999minI, comp2999minJ;
    Comparator comp2999(comp2272minVal, comp2272minI, comp2272minJ, comp2273minVal, comp2273minI, comp2273minJ, comp2999minVal, comp2999minI, comp2999minJ);
    wire [11:0] comp3000minVal;
    wire [5:0] comp3000minI, comp3000minJ;
    Comparator comp3000(comp2274minVal, comp2274minI, comp2274minJ, comp2275minVal, comp2275minI, comp2275minJ, comp3000minVal, comp3000minI, comp3000minJ);
    wire [11:0] comp3001minVal;
    wire [5:0] comp3001minI, comp3001minJ;
    Comparator comp3001(comp2276minVal, comp2276minI, comp2276minJ, comp2277minVal, comp2277minI, comp2277minJ, comp3001minVal, comp3001minI, comp3001minJ);
    wire [11:0] comp3002minVal;
    wire [5:0] comp3002minI, comp3002minJ;
    Comparator comp3002(comp2278minVal, comp2278minI, comp2278minJ, comp2279minVal, comp2279minI, comp2279minJ, comp3002minVal, comp3002minI, comp3002minJ);
    wire [11:0] comp3003minVal;
    wire [5:0] comp3003minI, comp3003minJ;
    Comparator comp3003(comp2280minVal, comp2280minI, comp2280minJ, comp2281minVal, comp2281minI, comp2281minJ, comp3003minVal, comp3003minI, comp3003minJ);
    wire [11:0] comp3004minVal;
    wire [5:0] comp3004minI, comp3004minJ;
    Comparator comp3004(comp2282minVal, comp2282minI, comp2282minJ, comp2283minVal, comp2283minI, comp2283minJ, comp3004minVal, comp3004minI, comp3004minJ);
    wire [11:0] comp3005minVal;
    wire [5:0] comp3005minI, comp3005minJ;
    Comparator comp3005(comp2284minVal, comp2284minI, comp2284minJ, comp2285minVal, comp2285minI, comp2285minJ, comp3005minVal, comp3005minI, comp3005minJ);
    wire [11:0] comp3006minVal;
    wire [5:0] comp3006minI, comp3006minJ;
    Comparator comp3006(comp2286minVal, comp2286minI, comp2286minJ, comp2287minVal, comp2287minI, comp2287minJ, comp3006minVal, comp3006minI, comp3006minJ);
    wire [11:0] comp3007minVal;
    wire [5:0] comp3007minI, comp3007minJ;
    Comparator comp3007(comp2288minVal, comp2288minI, comp2288minJ, comp2289minVal, comp2289minI, comp2289minJ, comp3007minVal, comp3007minI, comp3007minJ);
    wire [11:0] comp3008minVal;
    wire [5:0] comp3008minI, comp3008minJ;
    Comparator comp3008(comp2290minVal, comp2290minI, comp2290minJ, comp2291minVal, comp2291minI, comp2291minJ, comp3008minVal, comp3008minI, comp3008minJ);
    wire [11:0] comp3009minVal;
    wire [5:0] comp3009minI, comp3009minJ;
    Comparator comp3009(comp2292minVal, comp2292minI, comp2292minJ, comp2293minVal, comp2293minI, comp2293minJ, comp3009minVal, comp3009minI, comp3009minJ);
    wire [11:0] comp3010minVal;
    wire [5:0] comp3010minI, comp3010minJ;
    Comparator comp3010(comp2294minVal, comp2294minI, comp2294minJ, comp2295minVal, comp2295minI, comp2295minJ, comp3010minVal, comp3010minI, comp3010minJ);
    wire [11:0] comp3011minVal;
    wire [5:0] comp3011minI, comp3011minJ;
    Comparator comp3011(comp2296minVal, comp2296minI, comp2296minJ, comp2297minVal, comp2297minI, comp2297minJ, comp3011minVal, comp3011minI, comp3011minJ);
    wire [11:0] comp3012minVal;
    wire [5:0] comp3012minI, comp3012minJ;
    Comparator comp3012(comp2298minVal, comp2298minI, comp2298minJ, comp2299minVal, comp2299minI, comp2299minJ, comp3012minVal, comp3012minI, comp3012minJ);
    wire [11:0] comp3013minVal;
    wire [5:0] comp3013minI, comp3013minJ;
    Comparator comp3013(comp2300minVal, comp2300minI, comp2300minJ, comp2301minVal, comp2301minI, comp2301minJ, comp3013minVal, comp3013minI, comp3013minJ);
    wire [11:0] comp3014minVal;
    wire [5:0] comp3014minI, comp3014minJ;
    Comparator comp3014(comp2302minVal, comp2302minI, comp2302minJ, comp2303minVal, comp2303minI, comp2303minJ, comp3014minVal, comp3014minI, comp3014minJ);
    wire [11:0] comp3015minVal;
    wire [5:0] comp3015minI, comp3015minJ;
    Comparator comp3015(comp2304minVal, comp2304minI, comp2304minJ, comp2305minVal, comp2305minI, comp2305minJ, comp3015minVal, comp3015minI, comp3015minJ);
    wire [11:0] comp3016minVal;
    wire [5:0] comp3016minI, comp3016minJ;
    Comparator comp3016(comp2306minVal, comp2306minI, comp2306minJ, comp2307minVal, comp2307minI, comp2307minJ, comp3016minVal, comp3016minI, comp3016minJ);
    wire [11:0] comp3017minVal;
    wire [5:0] comp3017minI, comp3017minJ;
    Comparator comp3017(comp2308minVal, comp2308minI, comp2308minJ, comp2309minVal, comp2309minI, comp2309minJ, comp3017minVal, comp3017minI, comp3017minJ);
    wire [11:0] comp3018minVal;
    wire [5:0] comp3018minI, comp3018minJ;
    Comparator comp3018(comp2310minVal, comp2310minI, comp2310minJ, comp2311minVal, comp2311minI, comp2311minJ, comp3018minVal, comp3018minI, comp3018minJ);
    wire [11:0] comp3019minVal;
    wire [5:0] comp3019minI, comp3019minJ;
    Comparator comp3019(comp2312minVal, comp2312minI, comp2312minJ, comp2313minVal, comp2313minI, comp2313minJ, comp3019minVal, comp3019minI, comp3019minJ);
    wire [11:0] comp3020minVal;
    wire [5:0] comp3020minI, comp3020minJ;
    Comparator comp3020(comp2314minVal, comp2314minI, comp2314minJ, comp2315minVal, comp2315minI, comp2315minJ, comp3020minVal, comp3020minI, comp3020minJ);
    wire [11:0] comp3021minVal;
    wire [5:0] comp3021minI, comp3021minJ;
    Comparator comp3021(comp2316minVal, comp2316minI, comp2316minJ, comp2317minVal, comp2317minI, comp2317minJ, comp3021minVal, comp3021minI, comp3021minJ);
    wire [11:0] comp3022minVal;
    wire [5:0] comp3022minI, comp3022minJ;
    Comparator comp3022(comp2318minVal, comp2318minI, comp2318minJ, comp2319minVal, comp2319minI, comp2319minJ, comp3022minVal, comp3022minI, comp3022minJ);
    wire [11:0] comp3023minVal;
    wire [5:0] comp3023minI, comp3023minJ;
    Comparator comp3023(comp2320minVal, comp2320minI, comp2320minJ, comp2321minVal, comp2321minI, comp2321minJ, comp3023minVal, comp3023minI, comp3023minJ);
    wire [11:0] comp3024minVal;
    wire [5:0] comp3024minI, comp3024minJ;
    Comparator comp3024(comp2322minVal, comp2322minI, comp2322minJ, comp2323minVal, comp2323minI, comp2323minJ, comp3024minVal, comp3024minI, comp3024minJ);
    wire [11:0] comp3025minVal;
    wire [5:0] comp3025minI, comp3025minJ;
    Comparator comp3025(comp2324minVal, comp2324minI, comp2324minJ, comp2325minVal, comp2325minI, comp2325minJ, comp3025minVal, comp3025minI, comp3025minJ);
    wire [11:0] comp3026minVal;
    wire [5:0] comp3026minI, comp3026minJ;
    Comparator comp3026(comp2326minVal, comp2326minI, comp2326minJ, comp2327minVal, comp2327minI, comp2327minJ, comp3026minVal, comp3026minI, comp3026minJ);
    wire [11:0] comp3027minVal;
    wire [5:0] comp3027minI, comp3027minJ;
    Comparator comp3027(comp2328minVal, comp2328minI, comp2328minJ, comp2329minVal, comp2329minI, comp2329minJ, comp3027minVal, comp3027minI, comp3027minJ);
    wire [11:0] comp3028minVal;
    wire [5:0] comp3028minI, comp3028minJ;
    Comparator comp3028(comp2330minVal, comp2330minI, comp2330minJ, comp2331minVal, comp2331minI, comp2331minJ, comp3028minVal, comp3028minI, comp3028minJ);
    wire [11:0] comp3029minVal;
    wire [5:0] comp3029minI, comp3029minJ;
    Comparator comp3029(comp2332minVal, comp2332minI, comp2332minJ, comp2333minVal, comp2333minI, comp2333minJ, comp3029minVal, comp3029minI, comp3029minJ);
    wire [11:0] comp3030minVal;
    wire [5:0] comp3030minI, comp3030minJ;
    Comparator comp3030(comp2334minVal, comp2334minI, comp2334minJ, comp2335minVal, comp2335minI, comp2335minJ, comp3030minVal, comp3030minI, comp3030minJ);
    wire [11:0] comp3031minVal;
    wire [5:0] comp3031minI, comp3031minJ;
    Comparator comp3031(comp2336minVal, comp2336minI, comp2336minJ, comp2337minVal, comp2337minI, comp2337minJ, comp3031minVal, comp3031minI, comp3031minJ);
    wire [11:0] comp3032minVal;
    wire [5:0] comp3032minI, comp3032minJ;
    Comparator comp3032(comp2338minVal, comp2338minI, comp2338minJ, comp2339minVal, comp2339minI, comp2339minJ, comp3032minVal, comp3032minI, comp3032minJ);
    wire [11:0] comp3033minVal;
    wire [5:0] comp3033minI, comp3033minJ;
    Comparator comp3033(comp2340minVal, comp2340minI, comp2340minJ, comp2341minVal, comp2341minI, comp2341minJ, comp3033minVal, comp3033minI, comp3033minJ);
    wire [11:0] comp3034minVal;
    wire [5:0] comp3034minI, comp3034minJ;
    Comparator comp3034(comp2342minVal, comp2342minI, comp2342minJ, comp2343minVal, comp2343minI, comp2343minJ, comp3034minVal, comp3034minI, comp3034minJ);
    wire [11:0] comp3035minVal;
    wire [5:0] comp3035minI, comp3035minJ;
    Comparator comp3035(comp2344minVal, comp2344minI, comp2344minJ, comp2345minVal, comp2345minI, comp2345minJ, comp3035minVal, comp3035minI, comp3035minJ);
    wire [11:0] comp3036minVal;
    wire [5:0] comp3036minI, comp3036minJ;
    Comparator comp3036(comp2346minVal, comp2346minI, comp2346minJ, comp2347minVal, comp2347minI, comp2347minJ, comp3036minVal, comp3036minI, comp3036minJ);
    wire [11:0] comp3037minVal;
    wire [5:0] comp3037minI, comp3037minJ;
    Comparator comp3037(comp2348minVal, comp2348minI, comp2348minJ, comp2349minVal, comp2349minI, comp2349minJ, comp3037minVal, comp3037minI, comp3037minJ);
    wire [11:0] comp3038minVal;
    wire [5:0] comp3038minI, comp3038minJ;
    Comparator comp3038(comp2350minVal, comp2350minI, comp2350minJ, comp2351minVal, comp2351minI, comp2351minJ, comp3038minVal, comp3038minI, comp3038minJ);
    wire [11:0] comp3039minVal;
    wire [5:0] comp3039minI, comp3039minJ;
    Comparator comp3039(comp2352minVal, comp2352minI, comp2352minJ, comp2353minVal, comp2353minI, comp2353minJ, comp3039minVal, comp3039minI, comp3039minJ);
    wire [11:0] comp3040minVal;
    wire [5:0] comp3040minI, comp3040minJ;
    Comparator comp3040(comp2354minVal, comp2354minI, comp2354minJ, comp2355minVal, comp2355minI, comp2355minJ, comp3040minVal, comp3040minI, comp3040minJ);
    wire [11:0] comp3041minVal;
    wire [5:0] comp3041minI, comp3041minJ;
    Comparator comp3041(comp2356minVal, comp2356minI, comp2356minJ, comp2357minVal, comp2357minI, comp2357minJ, comp3041minVal, comp3041minI, comp3041minJ);
    wire [11:0] comp3042minVal;
    wire [5:0] comp3042minI, comp3042minJ;
    Comparator comp3042(comp2358minVal, comp2358minI, comp2358minJ, comp2359minVal, comp2359minI, comp2359minJ, comp3042minVal, comp3042minI, comp3042minJ);
    wire [11:0] comp3043minVal;
    wire [5:0] comp3043minI, comp3043minJ;
    Comparator comp3043(comp2360minVal, comp2360minI, comp2360minJ, comp2361minVal, comp2361minI, comp2361minJ, comp3043minVal, comp3043minI, comp3043minJ);
    wire [11:0] comp3044minVal;
    wire [5:0] comp3044minI, comp3044minJ;
    Comparator comp3044(comp2362minVal, comp2362minI, comp2362minJ, comp2363minVal, comp2363minI, comp2363minJ, comp3044minVal, comp3044minI, comp3044minJ);
    wire [11:0] comp3045minVal;
    wire [5:0] comp3045minI, comp3045minJ;
    Comparator comp3045(comp2364minVal, comp2364minI, comp2364minJ, comp2365minVal, comp2365minI, comp2365minJ, comp3045minVal, comp3045minI, comp3045minJ);
    wire [11:0] comp3046minVal;
    wire [5:0] comp3046minI, comp3046minJ;
    Comparator comp3046(comp2366minVal, comp2366minI, comp2366minJ, comp2367minVal, comp2367minI, comp2367minJ, comp3046minVal, comp3046minI, comp3046minJ);
    wire [11:0] comp3047minVal;
    wire [5:0] comp3047minI, comp3047minJ;
    Comparator comp3047(comp2368minVal, comp2368minI, comp2368minJ, comp2369minVal, comp2369minI, comp2369minJ, comp3047minVal, comp3047minI, comp3047minJ);
    wire [11:0] comp3048minVal;
    wire [5:0] comp3048minI, comp3048minJ;
    Comparator comp3048(comp2370minVal, comp2370minI, comp2370minJ, comp2371minVal, comp2371minI, comp2371minJ, comp3048minVal, comp3048minI, comp3048minJ);
    wire [11:0] comp3049minVal;
    wire [5:0] comp3049minI, comp3049minJ;
    Comparator comp3049(comp2372minVal, comp2372minI, comp2372minJ, comp2373minVal, comp2373minI, comp2373minJ, comp3049minVal, comp3049minI, comp3049minJ);
    wire [11:0] comp3050minVal;
    wire [5:0] comp3050minI, comp3050minJ;
    Comparator comp3050(comp2374minVal, comp2374minI, comp2374minJ, comp2375minVal, comp2375minI, comp2375minJ, comp3050minVal, comp3050minI, comp3050minJ);
    wire [11:0] comp3051minVal;
    wire [5:0] comp3051minI, comp3051minJ;
    Comparator comp3051(comp2376minVal, comp2376minI, comp2376minJ, comp2377minVal, comp2377minI, comp2377minJ, comp3051minVal, comp3051minI, comp3051minJ);
    wire [11:0] comp3052minVal;
    wire [5:0] comp3052minI, comp3052minJ;
    Comparator comp3052(comp2378minVal, comp2378minI, comp2378minJ, comp2379minVal, comp2379minI, comp2379minJ, comp3052minVal, comp3052minI, comp3052minJ);
    wire [11:0] comp3053minVal;
    wire [5:0] comp3053minI, comp3053minJ;
    Comparator comp3053(comp2380minVal, comp2380minI, comp2380minJ, comp2381minVal, comp2381minI, comp2381minJ, comp3053minVal, comp3053minI, comp3053minJ);
    wire [11:0] comp3054minVal;
    wire [5:0] comp3054minI, comp3054minJ;
    Comparator comp3054(comp2382minVal, comp2382minI, comp2382minJ, comp2383minVal, comp2383minI, comp2383minJ, comp3054minVal, comp3054minI, comp3054minJ);
    wire [11:0] comp3055minVal;
    wire [5:0] comp3055minI, comp3055minJ;
    Comparator comp3055(comp2384minVal, comp2384minI, comp2384minJ, comp2385minVal, comp2385minI, comp2385minJ, comp3055minVal, comp3055minI, comp3055minJ);
    wire [11:0] comp3056minVal;
    wire [5:0] comp3056minI, comp3056minJ;
    Comparator comp3056(comp2386minVal, comp2386minI, comp2386minJ, comp2387minVal, comp2387minI, comp2387minJ, comp3056minVal, comp3056minI, comp3056minJ);
    wire [11:0] comp3057minVal;
    wire [5:0] comp3057minI, comp3057minJ;
    Comparator comp3057(comp2388minVal, comp2388minI, comp2388minJ, comp2389minVal, comp2389minI, comp2389minJ, comp3057minVal, comp3057minI, comp3057minJ);
    wire [11:0] comp3058minVal;
    wire [5:0] comp3058minI, comp3058minJ;
    Comparator comp3058(comp2390minVal, comp2390minI, comp2390minJ, comp2391minVal, comp2391minI, comp2391minJ, comp3058minVal, comp3058minI, comp3058minJ);
    wire [11:0] comp3059minVal;
    wire [5:0] comp3059minI, comp3059minJ;
    Comparator comp3059(comp2392minVal, comp2392minI, comp2392minJ, comp2393minVal, comp2393minI, comp2393minJ, comp3059minVal, comp3059minI, comp3059minJ);
    wire [11:0] comp3060minVal;
    wire [5:0] comp3060minI, comp3060minJ;
    Comparator comp3060(comp2394minVal, comp2394minI, comp2394minJ, comp2395minVal, comp2395minI, comp2395minJ, comp3060minVal, comp3060minI, comp3060minJ);
    wire [11:0] comp3061minVal;
    wire [5:0] comp3061minI, comp3061minJ;
    Comparator comp3061(comp2396minVal, comp2396minI, comp2396minJ, comp2397minVal, comp2397minI, comp2397minJ, comp3061minVal, comp3061minI, comp3061minJ);
    wire [11:0] comp3062minVal;
    wire [5:0] comp3062minI, comp3062minJ;
    Comparator comp3062(comp2398minVal, comp2398minI, comp2398minJ, comp2399minVal, comp2399minI, comp2399minJ, comp3062minVal, comp3062minI, comp3062minJ);
    wire [11:0] comp3063minVal;
    wire [5:0] comp3063minI, comp3063minJ;
    Comparator comp3063(comp2400minVal, comp2400minI, comp2400minJ, comp2401minVal, comp2401minI, comp2401minJ, comp3063minVal, comp3063minI, comp3063minJ);
    wire [11:0] comp3064minVal;
    wire [5:0] comp3064minI, comp3064minJ;
    Comparator comp3064(comp2402minVal, comp2402minI, comp2402minJ, comp2403minVal, comp2403minI, comp2403minJ, comp3064minVal, comp3064minI, comp3064minJ);
    wire [11:0] comp3065minVal;
    wire [5:0] comp3065minI, comp3065minJ;
    Comparator comp3065(comp2404minVal, comp2404minI, comp2404minJ, comp2405minVal, comp2405minI, comp2405minJ, comp3065minVal, comp3065minI, comp3065minJ);
    wire [11:0] comp3066minVal;
    wire [5:0] comp3066minI, comp3066minJ;
    Comparator comp3066(comp2406minVal, comp2406minI, comp2406minJ, comp2407minVal, comp2407minI, comp2407minJ, comp3066minVal, comp3066minI, comp3066minJ);
    wire [11:0] comp3067minVal;
    wire [5:0] comp3067minI, comp3067minJ;
    Comparator comp3067(comp2408minVal, comp2408minI, comp2408minJ, comp2409minVal, comp2409minI, comp2409minJ, comp3067minVal, comp3067minI, comp3067minJ);
    wire [11:0] comp3068minVal;
    wire [5:0] comp3068minI, comp3068minJ;
    Comparator comp3068(comp2410minVal, comp2410minI, comp2410minJ, comp2411minVal, comp2411minI, comp2411minJ, comp3068minVal, comp3068minI, comp3068minJ);
    wire [11:0] comp3069minVal;
    wire [5:0] comp3069minI, comp3069minJ;
    Comparator comp3069(comp2412minVal, comp2412minI, comp2412minJ, comp2413minVal, comp2413minI, comp2413minJ, comp3069minVal, comp3069minI, comp3069minJ);
    wire [11:0] comp3070minVal;
    wire [5:0] comp3070minI, comp3070minJ;
    Comparator comp3070(comp2414minVal, comp2414minI, comp2414minJ, comp2415minVal, comp2415minI, comp2415minJ, comp3070minVal, comp3070minI, comp3070minJ);
    wire [11:0] comp3071minVal;
    wire [5:0] comp3071minI, comp3071minJ;
    Comparator comp3071(comp2416minVal, comp2416minI, comp2416minJ, comp2417minVal, comp2417minI, comp2417minJ, comp3071minVal, comp3071minI, comp3071minJ);
    wire [11:0] comp3072minVal;
    wire [5:0] comp3072minI, comp3072minJ;
    Comparator comp3072(comp2418minVal, comp2418minI, comp2418minJ, comp2419minVal, comp2419minI, comp2419minJ, comp3072minVal, comp3072minI, comp3072minJ);
    wire [11:0] comp3073minVal;
    wire [5:0] comp3073minI, comp3073minJ;
    Comparator comp3073(comp2420minVal, comp2420minI, comp2420minJ, comp2421minVal, comp2421minI, comp2421minJ, comp3073minVal, comp3073minI, comp3073minJ);
    wire [11:0] comp3074minVal;
    wire [5:0] comp3074minI, comp3074minJ;
    Comparator comp3074(comp2422minVal, comp2422minI, comp2422minJ, comp2423minVal, comp2423minI, comp2423minJ, comp3074minVal, comp3074minI, comp3074minJ);
    wire [11:0] comp3075minVal;
    wire [5:0] comp3075minI, comp3075minJ;
    Comparator comp3075(comp2424minVal, comp2424minI, comp2424minJ, comp2425minVal, comp2425minI, comp2425minJ, comp3075minVal, comp3075minI, comp3075minJ);
    wire [11:0] comp3076minVal;
    wire [5:0] comp3076minI, comp3076minJ;
    Comparator comp3076(comp2426minVal, comp2426minI, comp2426minJ, comp2427minVal, comp2427minI, comp2427minJ, comp3076minVal, comp3076minI, comp3076minJ);
    wire [11:0] comp3077minVal;
    wire [5:0] comp3077minI, comp3077minJ;
    Comparator comp3077(comp2428minVal, comp2428minI, comp2428minJ, comp2429minVal, comp2429minI, comp2429minJ, comp3077minVal, comp3077minI, comp3077minJ);
    wire [11:0] comp3078minVal;
    wire [5:0] comp3078minI, comp3078minJ;
    Comparator comp3078(comp2430minVal, comp2430minI, comp2430minJ, comp2431minVal, comp2431minI, comp2431minJ, comp3078minVal, comp3078minI, comp3078minJ);
    wire [11:0] comp3079minVal;
    wire [5:0] comp3079minI, comp3079minJ;
    Comparator comp3079(comp2432minVal, comp2432minI, comp2432minJ, comp2433minVal, comp2433minI, comp2433minJ, comp3079minVal, comp3079minI, comp3079minJ);
    wire [11:0] comp3080minVal;
    wire [5:0] comp3080minI, comp3080minJ;
    Comparator comp3080(comp2434minVal, comp2434minI, comp2434minJ, comp2435minVal, comp2435minI, comp2435minJ, comp3080minVal, comp3080minI, comp3080minJ);
    wire [11:0] comp3081minVal;
    wire [5:0] comp3081minI, comp3081minJ;
    Comparator comp3081(comp2436minVal, comp2436minI, comp2436minJ, comp2437minVal, comp2437minI, comp2437minJ, comp3081minVal, comp3081minI, comp3081minJ);
    wire [11:0] comp3082minVal;
    wire [5:0] comp3082minI, comp3082minJ;
    Comparator comp3082(comp2438minVal, comp2438minI, comp2438minJ, comp2439minVal, comp2439minI, comp2439minJ, comp3082minVal, comp3082minI, comp3082minJ);
    wire [11:0] comp3083minVal;
    wire [5:0] comp3083minI, comp3083minJ;
    Comparator comp3083(comp2440minVal, comp2440minI, comp2440minJ, comp2441minVal, comp2441minI, comp2441minJ, comp3083minVal, comp3083minI, comp3083minJ);
    wire [11:0] comp3084minVal;
    wire [5:0] comp3084minI, comp3084minJ;
    Comparator comp3084(comp2442minVal, comp2442minI, comp2442minJ, comp2443minVal, comp2443minI, comp2443minJ, comp3084minVal, comp3084minI, comp3084minJ);
    wire [11:0] comp3085minVal;
    wire [5:0] comp3085minI, comp3085minJ;
    Comparator comp3085(comp2444minVal, comp2444minI, comp2444minJ, comp2445minVal, comp2445minI, comp2445minJ, comp3085minVal, comp3085minI, comp3085minJ);
    wire [11:0] comp3086minVal;
    wire [5:0] comp3086minI, comp3086minJ;
    Comparator comp3086(comp2446minVal, comp2446minI, comp2446minJ, comp2447minVal, comp2447minI, comp2447minJ, comp3086minVal, comp3086minI, comp3086minJ);
    wire [11:0] comp3087minVal;
    wire [5:0] comp3087minI, comp3087minJ;
    Comparator comp3087(comp2448minVal, comp2448minI, comp2448minJ, comp2449minVal, comp2449minI, comp2449minJ, comp3087minVal, comp3087minI, comp3087minJ);
    wire [11:0] comp3088minVal;
    wire [5:0] comp3088minI, comp3088minJ;
    Comparator comp3088(comp2450minVal, comp2450minI, comp2450minJ, comp2451minVal, comp2451minI, comp2451minJ, comp3088minVal, comp3088minI, comp3088minJ);
    wire [11:0] comp3089minVal;
    wire [5:0] comp3089minI, comp3089minJ;
    Comparator comp3089(comp2452minVal, comp2452minI, comp2452minJ, comp2453minVal, comp2453minI, comp2453minJ, comp3089minVal, comp3089minI, comp3089minJ);
    wire [11:0] comp3090minVal;
    wire [5:0] comp3090minI, comp3090minJ;
    Comparator comp3090(comp2454minVal, comp2454minI, comp2454minJ, comp2455minVal, comp2455minI, comp2455minJ, comp3090minVal, comp3090minI, comp3090minJ);
    wire [11:0] comp3091minVal;
    wire [5:0] comp3091minI, comp3091minJ;
    Comparator comp3091(comp2456minVal, comp2456minI, comp2456minJ, comp2457minVal, comp2457minI, comp2457minJ, comp3091minVal, comp3091minI, comp3091minJ);
    wire [11:0] comp3092minVal;
    wire [5:0] comp3092minI, comp3092minJ;
    Comparator comp3092(comp2458minVal, comp2458minI, comp2458minJ, comp2459minVal, comp2459minI, comp2459minJ, comp3092minVal, comp3092minI, comp3092minJ);
    wire [11:0] comp3093minVal;
    wire [5:0] comp3093minI, comp3093minJ;
    Comparator comp3093(comp2460minVal, comp2460minI, comp2460minJ, comp2461minVal, comp2461minI, comp2461minJ, comp3093minVal, comp3093minI, comp3093minJ);
    wire [11:0] comp3094minVal;
    wire [5:0] comp3094minI, comp3094minJ;
    Comparator comp3094(comp2462minVal, comp2462minI, comp2462minJ, comp2463minVal, comp2463minI, comp2463minJ, comp3094minVal, comp3094minI, comp3094minJ);
    wire [11:0] comp3095minVal;
    wire [5:0] comp3095minI, comp3095minJ;
    Comparator comp3095(comp2464minVal, comp2464minI, comp2464minJ, comp2465minVal, comp2465minI, comp2465minJ, comp3095minVal, comp3095minI, comp3095minJ);
    wire [11:0] comp3096minVal;
    wire [5:0] comp3096minI, comp3096minJ;
    Comparator comp3096(comp2466minVal, comp2466minI, comp2466minJ, comp2467minVal, comp2467minI, comp2467minJ, comp3096minVal, comp3096minI, comp3096minJ);
    wire [11:0] comp3097minVal;
    wire [5:0] comp3097minI, comp3097minJ;
    Comparator comp3097(comp2468minVal, comp2468minI, comp2468minJ, comp2469minVal, comp2469minI, comp2469minJ, comp3097minVal, comp3097minI, comp3097minJ);
    wire [11:0] comp3098minVal;
    wire [5:0] comp3098minI, comp3098minJ;
    Comparator comp3098(comp2470minVal, comp2470minI, comp2470minJ, comp2471minVal, comp2471minI, comp2471minJ, comp3098minVal, comp3098minI, comp3098minJ);
    wire [11:0] comp3099minVal;
    wire [5:0] comp3099minI, comp3099minJ;
    Comparator comp3099(comp2472minVal, comp2472minI, comp2472minJ, comp2473minVal, comp2473minI, comp2473minJ, comp3099minVal, comp3099minI, comp3099minJ);
    wire [11:0] comp3100minVal;
    wire [5:0] comp3100minI, comp3100minJ;
    Comparator comp3100(comp2474minVal, comp2474minI, comp2474minJ, comp2475minVal, comp2475minI, comp2475minJ, comp3100minVal, comp3100minI, comp3100minJ);
    wire [11:0] comp3101minVal;
    wire [5:0] comp3101minI, comp3101minJ;
    Comparator comp3101(comp2476minVal, comp2476minI, comp2476minJ, comp2477minVal, comp2477minI, comp2477minJ, comp3101minVal, comp3101minI, comp3101minJ);
    wire [11:0] comp3102minVal;
    wire [5:0] comp3102minI, comp3102minJ;
    Comparator comp3102(comp2478minVal, comp2478minI, comp2478minJ, comp2479minVal, comp2479minI, comp2479minJ, comp3102minVal, comp3102minI, comp3102minJ);
    wire [11:0] comp3103minVal;
    wire [5:0] comp3103minI, comp3103minJ;
    Comparator comp3103(comp2480minVal, comp2480minI, comp2480minJ, comp2481minVal, comp2481minI, comp2481minJ, comp3103minVal, comp3103minI, comp3103minJ);
    wire [11:0] comp3104minVal;
    wire [5:0] comp3104minI, comp3104minJ;
    Comparator comp3104(comp2482minVal, comp2482minI, comp2482minJ, comp2483minVal, comp2483minI, comp2483minJ, comp3104minVal, comp3104minI, comp3104minJ);
    wire [11:0] comp3105minVal;
    wire [5:0] comp3105minI, comp3105minJ;
    Comparator comp3105(comp2484minVal, comp2484minI, comp2484minJ, comp2485minVal, comp2485minI, comp2485minJ, comp3105minVal, comp3105minI, comp3105minJ);
    wire [11:0] comp3106minVal;
    wire [5:0] comp3106minI, comp3106minJ;
    Comparator comp3106(comp2486minVal, comp2486minI, comp2486minJ, comp2487minVal, comp2487minI, comp2487minJ, comp3106minVal, comp3106minI, comp3106minJ);
    wire [11:0] comp3107minVal;
    wire [5:0] comp3107minI, comp3107minJ;
    Comparator comp3107(comp2488minVal, comp2488minI, comp2488minJ, comp2489minVal, comp2489minI, comp2489minJ, comp3107minVal, comp3107minI, comp3107minJ);
    wire [11:0] comp3108minVal;
    wire [5:0] comp3108minI, comp3108minJ;
    Comparator comp3108(comp2490minVal, comp2490minI, comp2490minJ, comp2491minVal, comp2491minI, comp2491minJ, comp3108minVal, comp3108minI, comp3108minJ);
    wire [11:0] comp3109minVal;
    wire [5:0] comp3109minI, comp3109minJ;
    Comparator comp3109(comp2492minVal, comp2492minI, comp2492minJ, comp2493minVal, comp2493minI, comp2493minJ, comp3109minVal, comp3109minI, comp3109minJ);
    wire [11:0] comp3110minVal;
    wire [5:0] comp3110minI, comp3110minJ;
    Comparator comp3110(comp2494minVal, comp2494minI, comp2494minJ, comp2495minVal, comp2495minI, comp2495minJ, comp3110minVal, comp3110minI, comp3110minJ);
    wire [11:0] comp3111minVal;
    wire [5:0] comp3111minI, comp3111minJ;
    Comparator comp3111(comp2496minVal, comp2496minI, comp2496minJ, comp2497minVal, comp2497minI, comp2497minJ, comp3111minVal, comp3111minI, comp3111minJ);
    wire [11:0] comp3112minVal;
    wire [5:0] comp3112minI, comp3112minJ;
    Comparator comp3112(comp2498minVal, comp2498minI, comp2498minJ, comp2499minVal, comp2499minI, comp2499minJ, comp3112minVal, comp3112minI, comp3112minJ);
    wire [11:0] comp3113minVal;
    wire [5:0] comp3113minI, comp3113minJ;
    Comparator comp3113(comp2500minVal, comp2500minI, comp2500minJ, comp2501minVal, comp2501minI, comp2501minJ, comp3113minVal, comp3113minI, comp3113minJ);
    wire [11:0] comp3114minVal;
    wire [5:0] comp3114minI, comp3114minJ;
    Comparator comp3114(comp2502minVal, comp2502minI, comp2502minJ, comp2503minVal, comp2503minI, comp2503minJ, comp3114minVal, comp3114minI, comp3114minJ);
    wire [11:0] comp3115minVal;
    wire [5:0] comp3115minI, comp3115minJ;
    Comparator comp3115(comp2504minVal, comp2504minI, comp2504minJ, comp2505minVal, comp2505minI, comp2505minJ, comp3115minVal, comp3115minI, comp3115minJ);
    wire [11:0] comp3116minVal;
    wire [5:0] comp3116minI, comp3116minJ;
    Comparator comp3116(comp2506minVal, comp2506minI, comp2506minJ, comp2507minVal, comp2507minI, comp2507minJ, comp3116minVal, comp3116minI, comp3116minJ);
    wire [11:0] comp3117minVal;
    wire [5:0] comp3117minI, comp3117minJ;
    Comparator comp3117(comp2508minVal, comp2508minI, comp2508minJ, comp2509minVal, comp2509minI, comp2509minJ, comp3117minVal, comp3117minI, comp3117minJ);
    wire [11:0] comp3118minVal;
    wire [5:0] comp3118minI, comp3118minJ;
    Comparator comp3118(comp2510minVal, comp2510minI, comp2510minJ, comp2511minVal, comp2511minI, comp2511minJ, comp3118minVal, comp3118minI, comp3118minJ);
    wire [11:0] comp3119minVal;
    wire [5:0] comp3119minI, comp3119minJ;
    Comparator comp3119(comp2512minVal, comp2512minI, comp2512minJ, comp2513minVal, comp2513minI, comp2513minJ, comp3119minVal, comp3119minI, comp3119minJ);
    wire [11:0] comp3120minVal;
    wire [5:0] comp3120minI, comp3120minJ;
    Comparator comp3120(comp2514minVal, comp2514minI, comp2514minJ, comp2515minVal, comp2515minI, comp2515minJ, comp3120minVal, comp3120minI, comp3120minJ);
    wire [11:0] comp3121minVal;
    wire [5:0] comp3121minI, comp3121minJ;
    Comparator comp3121(comp2516minVal, comp2516minI, comp2516minJ, comp2517minVal, comp2517minI, comp2517minJ, comp3121minVal, comp3121minI, comp3121minJ);
    wire [11:0] comp3122minVal;
    wire [5:0] comp3122minI, comp3122minJ;
    Comparator comp3122(comp2518minVal, comp2518minI, comp2518minJ, comp2519minVal, comp2519minI, comp2519minJ, comp3122minVal, comp3122minI, comp3122minJ);
    wire [11:0] comp3123minVal;
    wire [5:0] comp3123minI, comp3123minJ;
    Comparator comp3123(comp2520minVal, comp2520minI, comp2520minJ, comp2521minVal, comp2521minI, comp2521minJ, comp3123minVal, comp3123minI, comp3123minJ);
    wire [11:0] comp3124minVal;
    wire [5:0] comp3124minI, comp3124minJ;
    Comparator comp3124(comp2522minVal, comp2522minI, comp2522minJ, comp2523minVal, comp2523minI, comp2523minJ, comp3124minVal, comp3124minI, comp3124minJ);
    wire [11:0] comp3125minVal;
    wire [5:0] comp3125minI, comp3125minJ;
    Comparator comp3125(comp2524minVal, comp2524minI, comp2524minJ, comp2525minVal, comp2525minI, comp2525minJ, comp3125minVal, comp3125minI, comp3125minJ);
    wire [11:0] comp3126minVal;
    wire [5:0] comp3126minI, comp3126minJ;
    Comparator comp3126(comp2526minVal, comp2526minI, comp2526minJ, comp2527minVal, comp2527minI, comp2527minJ, comp3126minVal, comp3126minI, comp3126minJ);
    wire [11:0] comp3127minVal;
    wire [5:0] comp3127minI, comp3127minJ;
    Comparator comp3127(comp2528minVal, comp2528minI, comp2528minJ, comp2529minVal, comp2529minI, comp2529minJ, comp3127minVal, comp3127minI, comp3127minJ);
    wire [11:0] comp3128minVal;
    wire [5:0] comp3128minI, comp3128minJ;
    Comparator comp3128(comp2530minVal, comp2530minI, comp2530minJ, comp2531minVal, comp2531minI, comp2531minJ, comp3128minVal, comp3128minI, comp3128minJ);
    wire [11:0] comp3129minVal;
    wire [5:0] comp3129minI, comp3129minJ;
    Comparator comp3129(comp2532minVal, comp2532minI, comp2532minJ, comp2533minVal, comp2533minI, comp2533minJ, comp3129minVal, comp3129minI, comp3129minJ);
    wire [11:0] comp3130minVal;
    wire [5:0] comp3130minI, comp3130minJ;
    Comparator comp3130(comp2534minVal, comp2534minI, comp2534minJ, comp2535minVal, comp2535minI, comp2535minJ, comp3130minVal, comp3130minI, comp3130minJ);
    wire [11:0] comp3131minVal;
    wire [5:0] comp3131minI, comp3131minJ;
    Comparator comp3131(comp2536minVal, comp2536minI, comp2536minJ, comp2537minVal, comp2537minI, comp2537minJ, comp3131minVal, comp3131minI, comp3131minJ);
    wire [11:0] comp3132minVal;
    wire [5:0] comp3132minI, comp3132minJ;
    Comparator comp3132(comp2538minVal, comp2538minI, comp2538minJ, comp2539minVal, comp2539minI, comp2539minJ, comp3132minVal, comp3132minI, comp3132minJ);
    wire [11:0] comp3133minVal;
    wire [5:0] comp3133minI, comp3133minJ;
    Comparator comp3133(comp2540minVal, comp2540minI, comp2540minJ, comp2541minVal, comp2541minI, comp2541minJ, comp3133minVal, comp3133minI, comp3133minJ);
    wire [11:0] comp3134minVal;
    wire [5:0] comp3134minI, comp3134minJ;
    Comparator comp3134(comp2542minVal, comp2542minI, comp2542minJ, comp2543minVal, comp2543minI, comp2543minJ, comp3134minVal, comp3134minI, comp3134minJ);
    wire [11:0] comp3135minVal;
    wire [5:0] comp3135minI, comp3135minJ;
    Comparator comp3135(comp2544minVal, comp2544minI, comp2544minJ, comp2545minVal, comp2545minI, comp2545minJ, comp3135minVal, comp3135minI, comp3135minJ);
    wire [11:0] comp3136minVal;
    wire [5:0] comp3136minI, comp3136minJ;
    Comparator comp3136(comp2546minVal, comp2546minI, comp2546minJ, comp2547minVal, comp2547minI, comp2547minJ, comp3136minVal, comp3136minI, comp3136minJ);
    wire [11:0] comp3137minVal;
    wire [5:0] comp3137minI, comp3137minJ;
    Comparator comp3137(comp2548minVal, comp2548minI, comp2548minJ, comp2549minVal, comp2549minI, comp2549minJ, comp3137minVal, comp3137minI, comp3137minJ);
    wire [11:0] comp3138minVal;
    wire [5:0] comp3138minI, comp3138minJ;
    Comparator comp3138(comp2550minVal, comp2550minI, comp2550minJ, comp2551minVal, comp2551minI, comp2551minJ, comp3138minVal, comp3138minI, comp3138minJ);
    wire [11:0] comp3139minVal;
    wire [5:0] comp3139minI, comp3139minJ;
    Comparator comp3139(comp2552minVal, comp2552minI, comp2552minJ, comp2553minVal, comp2553minI, comp2553minJ, comp3139minVal, comp3139minI, comp3139minJ);
    wire [11:0] comp3140minVal;
    wire [5:0] comp3140minI, comp3140minJ;
    Comparator comp3140(comp2554minVal, comp2554minI, comp2554minJ, comp2555minVal, comp2555minI, comp2555minJ, comp3140minVal, comp3140minI, comp3140minJ);
    wire [11:0] comp3141minVal;
    wire [5:0] comp3141minI, comp3141minJ;
    Comparator comp3141(comp2556minVal, comp2556minI, comp2556minJ, comp2557minVal, comp2557minI, comp2557minJ, comp3141minVal, comp3141minI, comp3141minJ);
    wire [11:0] comp3142minVal;
    wire [5:0] comp3142minI, comp3142minJ;
    Comparator comp3142(comp2558minVal, comp2558minI, comp2558minJ, comp2559minVal, comp2559minI, comp2559minJ, comp3142minVal, comp3142minI, comp3142minJ);
    wire [11:0] comp3143minVal;
    wire [5:0] comp3143minI, comp3143minJ;
    Comparator comp3143(comp2560minVal, comp2560minI, comp2560minJ, comp2561minVal, comp2561minI, comp2561minJ, comp3143minVal, comp3143minI, comp3143minJ);
    wire [11:0] comp3144minVal;
    wire [5:0] comp3144minI, comp3144minJ;
    Comparator comp3144(comp2562minVal, comp2562minI, comp2562minJ, comp2563minVal, comp2563minI, comp2563minJ, comp3144minVal, comp3144minI, comp3144minJ);
    wire [11:0] comp3145minVal;
    wire [5:0] comp3145minI, comp3145minJ;
    Comparator comp3145(comp2564minVal, comp2564minI, comp2564minJ, comp2565minVal, comp2565minI, comp2565minJ, comp3145minVal, comp3145minI, comp3145minJ);
    wire [11:0] comp3146minVal;
    wire [5:0] comp3146minI, comp3146minJ;
    Comparator comp3146(comp2566minVal, comp2566minI, comp2566minJ, comp2567minVal, comp2567minI, comp2567minJ, comp3146minVal, comp3146minI, comp3146minJ);
    wire [11:0] comp3147minVal;
    wire [5:0] comp3147minI, comp3147minJ;
    Comparator comp3147(comp2568minVal, comp2568minI, comp2568minJ, comp2569minVal, comp2569minI, comp2569minJ, comp3147minVal, comp3147minI, comp3147minJ);
    wire [11:0] comp3148minVal;
    wire [5:0] comp3148minI, comp3148minJ;
    Comparator comp3148(comp2570minVal, comp2570minI, comp2570minJ, comp2571minVal, comp2571minI, comp2571minJ, comp3148minVal, comp3148minI, comp3148minJ);
    wire [11:0] comp3149minVal;
    wire [5:0] comp3149minI, comp3149minJ;
    Comparator comp3149(comp2572minVal, comp2572minI, comp2572minJ, comp2573minVal, comp2573minI, comp2573minJ, comp3149minVal, comp3149minI, comp3149minJ);
    wire [11:0] comp3150minVal;
    wire [5:0] comp3150minI, comp3150minJ;
    Comparator comp3150(comp2574minVal, comp2574minI, comp2574minJ, comp2575minVal, comp2575minI, comp2575minJ, comp3150minVal, comp3150minI, comp3150minJ);
    wire [11:0] comp3151minVal;
    wire [5:0] comp3151minI, comp3151minJ;
    Comparator comp3151(comp2576minVal, comp2576minI, comp2576minJ, comp2577minVal, comp2577minI, comp2577minJ, comp3151minVal, comp3151minI, comp3151minJ);
    wire [11:0] comp3152minVal;
    wire [5:0] comp3152minI, comp3152minJ;
    Comparator comp3152(comp2578minVal, comp2578minI, comp2578minJ, comp2579minVal, comp2579minI, comp2579minJ, comp3152minVal, comp3152minI, comp3152minJ);
    wire [11:0] comp3153minVal;
    wire [5:0] comp3153minI, comp3153minJ;
    Comparator comp3153(comp2580minVal, comp2580minI, comp2580minJ, comp2581minVal, comp2581minI, comp2581minJ, comp3153minVal, comp3153minI, comp3153minJ);
    wire [11:0] comp3154minVal;
    wire [5:0] comp3154minI, comp3154minJ;
    Comparator comp3154(comp2582minVal, comp2582minI, comp2582minJ, comp2583minVal, comp2583minI, comp2583minJ, comp3154minVal, comp3154minI, comp3154minJ);
    wire [11:0] comp3155minVal;
    wire [5:0] comp3155minI, comp3155minJ;
    Comparator comp3155(comp2584minVal, comp2584minI, comp2584minJ, comp2585minVal, comp2585minI, comp2585minJ, comp3155minVal, comp3155minI, comp3155minJ);
    wire [11:0] comp3156minVal;
    wire [5:0] comp3156minI, comp3156minJ;
    Comparator comp3156(comp2586minVal, comp2586minI, comp2586minJ, comp2587minVal, comp2587minI, comp2587minJ, comp3156minVal, comp3156minI, comp3156minJ);
    wire [11:0] comp3157minVal;
    wire [5:0] comp3157minI, comp3157minJ;
    Comparator comp3157(comp2588minVal, comp2588minI, comp2588minJ, comp2589minVal, comp2589minI, comp2589minJ, comp3157minVal, comp3157minI, comp3157minJ);
    wire [11:0] comp3158minVal;
    wire [5:0] comp3158minI, comp3158minJ;
    Comparator comp3158(comp2590minVal, comp2590minI, comp2590minJ, comp2591minVal, comp2591minI, comp2591minJ, comp3158minVal, comp3158minI, comp3158minJ);
    wire [11:0] comp3159minVal;
    wire [5:0] comp3159minI, comp3159minJ;
    Comparator comp3159(comp2592minVal, comp2592minI, comp2592minJ, comp2593minVal, comp2593minI, comp2593minJ, comp3159minVal, comp3159minI, comp3159minJ);
    wire [11:0] comp3160minVal;
    wire [5:0] comp3160minI, comp3160minJ;
    Comparator comp3160(comp2594minVal, comp2594minI, comp2594minJ, comp2595minVal, comp2595minI, comp2595minJ, comp3160minVal, comp3160minI, comp3160minJ);
    wire [11:0] comp3161minVal;
    wire [5:0] comp3161minI, comp3161minJ;
    Comparator comp3161(comp2596minVal, comp2596minI, comp2596minJ, comp2597minVal, comp2597minI, comp2597minJ, comp3161minVal, comp3161minI, comp3161minJ);
    wire [11:0] comp3162minVal;
    wire [5:0] comp3162minI, comp3162minJ;
    Comparator comp3162(comp2598minVal, comp2598minI, comp2598minJ, comp2599minVal, comp2599minI, comp2599minJ, comp3162minVal, comp3162minI, comp3162minJ);
    wire [11:0] comp3163minVal;
    wire [5:0] comp3163minI, comp3163minJ;
    Comparator comp3163(comp2600minVal, comp2600minI, comp2600minJ, comp2601minVal, comp2601minI, comp2601minJ, comp3163minVal, comp3163minI, comp3163minJ);
    wire [11:0] comp3164minVal;
    wire [5:0] comp3164minI, comp3164minJ;
    Comparator comp3164(comp2602minVal, comp2602minI, comp2602minJ, comp2603minVal, comp2603minI, comp2603minJ, comp3164minVal, comp3164minI, comp3164minJ);
    wire [11:0] comp3165minVal;
    wire [5:0] comp3165minI, comp3165minJ;
    Comparator comp3165(comp2604minVal, comp2604minI, comp2604minJ, comp2605minVal, comp2605minI, comp2605minJ, comp3165minVal, comp3165minI, comp3165minJ);
    wire [11:0] comp3166minVal;
    wire [5:0] comp3166minI, comp3166minJ;
    Comparator comp3166(comp2606minVal, comp2606minI, comp2606minJ, comp2607minVal, comp2607minI, comp2607minJ, comp3166minVal, comp3166minI, comp3166minJ);
    wire [11:0] comp3167minVal;
    wire [5:0] comp3167minI, comp3167minJ;
    Comparator comp3167(comp2608minVal, comp2608minI, comp2608minJ, comp2609minVal, comp2609minI, comp2609minJ, comp3167minVal, comp3167minI, comp3167minJ);
    wire [11:0] comp3168minVal;
    wire [5:0] comp3168minI, comp3168minJ;
    Comparator comp3168(comp2610minVal, comp2610minI, comp2610minJ, comp2611minVal, comp2611minI, comp2611minJ, comp3168minVal, comp3168minI, comp3168minJ);
    wire [11:0] comp3169minVal;
    wire [5:0] comp3169minI, comp3169minJ;
    Comparator comp3169(comp2612minVal, comp2612minI, comp2612minJ, comp2613minVal, comp2613minI, comp2613minJ, comp3169minVal, comp3169minI, comp3169minJ);
    wire [11:0] comp3170minVal;
    wire [5:0] comp3170minI, comp3170minJ;
    Comparator comp3170(comp2614minVal, comp2614minI, comp2614minJ, comp2615minVal, comp2615minI, comp2615minJ, comp3170minVal, comp3170minI, comp3170minJ);
    wire [11:0] comp3171minVal;
    wire [5:0] comp3171minI, comp3171minJ;
    Comparator comp3171(comp2616minVal, comp2616minI, comp2616minJ, comp2617minVal, comp2617minI, comp2617minJ, comp3171minVal, comp3171minI, comp3171minJ);
    wire [11:0] comp3172minVal;
    wire [5:0] comp3172minI, comp3172minJ;
    Comparator comp3172(comp2618minVal, comp2618minI, comp2618minJ, comp2619minVal, comp2619minI, comp2619minJ, comp3172minVal, comp3172minI, comp3172minJ);
    wire [11:0] comp3173minVal;
    wire [5:0] comp3173minI, comp3173minJ;
    Comparator comp3173(comp2620minVal, comp2620minI, comp2620minJ, comp2621minVal, comp2621minI, comp2621minJ, comp3173minVal, comp3173minI, comp3173minJ);
    wire [11:0] comp3174minVal;
    wire [5:0] comp3174minI, comp3174minJ;
    Comparator comp3174(comp2622minVal, comp2622minI, comp2622minJ, comp2623minVal, comp2623minI, comp2623minJ, comp3174minVal, comp3174minI, comp3174minJ);
    wire [11:0] comp3175minVal;
    wire [5:0] comp3175minI, comp3175minJ;
    Comparator comp3175(comp2624minVal, comp2624minI, comp2624minJ, comp2625minVal, comp2625minI, comp2625minJ, comp3175minVal, comp3175minI, comp3175minJ);
    wire [11:0] comp3176minVal;
    wire [5:0] comp3176minI, comp3176minJ;
    Comparator comp3176(comp2626minVal, comp2626minI, comp2626minJ, comp2627minVal, comp2627minI, comp2627minJ, comp3176minVal, comp3176minI, comp3176minJ);
    wire [11:0] comp3177minVal;
    wire [5:0] comp3177minI, comp3177minJ;
    Comparator comp3177(comp2628minVal, comp2628minI, comp2628minJ, comp2629minVal, comp2629minI, comp2629minJ, comp3177minVal, comp3177minI, comp3177minJ);
    wire [11:0] comp3178minVal;
    wire [5:0] comp3178minI, comp3178minJ;
    Comparator comp3178(comp2630minVal, comp2630minI, comp2630minJ, comp2631minVal, comp2631minI, comp2631minJ, comp3178minVal, comp3178minI, comp3178minJ);
    wire [11:0] comp3179minVal;
    wire [5:0] comp3179minI, comp3179minJ;
    Comparator comp3179(comp2632minVal, comp2632minI, comp2632minJ, comp2633minVal, comp2633minI, comp2633minJ, comp3179minVal, comp3179minI, comp3179minJ);
    wire [11:0] comp3180minVal;
    wire [5:0] comp3180minI, comp3180minJ;
    Comparator comp3180(comp2634minVal, comp2634minI, comp2634minJ, comp2635minVal, comp2635minI, comp2635minJ, comp3180minVal, comp3180minI, comp3180minJ);
    wire [11:0] comp3181minVal;
    wire [5:0] comp3181minI, comp3181minJ;
    Comparator comp3181(comp2636minVal, comp2636minI, comp2636minJ, comp2637minVal, comp2637minI, comp2637minJ, comp3181minVal, comp3181minI, comp3181minJ);
    wire [11:0] comp3182minVal;
    wire [5:0] comp3182minI, comp3182minJ;
    Comparator comp3182(comp2638minVal, comp2638minI, comp2638minJ, comp2639minVal, comp2639minI, comp2639minJ, comp3182minVal, comp3182minI, comp3182minJ);
    wire [11:0] comp3183minVal;
    wire [5:0] comp3183minI, comp3183minJ;
    Comparator comp3183(comp2640minVal, comp2640minI, comp2640minJ, comp2641minVal, comp2641minI, comp2641minJ, comp3183minVal, comp3183minI, comp3183minJ);
    wire [11:0] comp3184minVal;
    wire [5:0] comp3184minI, comp3184minJ;
    Comparator comp3184(comp2642minVal, comp2642minI, comp2642minJ, comp2643minVal, comp2643minI, comp2643minJ, comp3184minVal, comp3184minI, comp3184minJ);
    wire [11:0] comp3185minVal;
    wire [5:0] comp3185minI, comp3185minJ;
    Comparator comp3185(comp2644minVal, comp2644minI, comp2644minJ, comp2645minVal, comp2645minI, comp2645minJ, comp3185minVal, comp3185minI, comp3185minJ);
    wire [11:0] comp3186minVal;
    wire [5:0] comp3186minI, comp3186minJ;
    Comparator comp3186(comp2646minVal, comp2646minI, comp2646minJ, comp2647minVal, comp2647minI, comp2647minJ, comp3186minVal, comp3186minI, comp3186minJ);
    wire [11:0] comp3187minVal;
    wire [5:0] comp3187minI, comp3187minJ;
    Comparator comp3187(comp2648minVal, comp2648minI, comp2648minJ, comp2649minVal, comp2649minI, comp2649minJ, comp3187minVal, comp3187minI, comp3187minJ);
    wire [11:0] comp3188minVal;
    wire [5:0] comp3188minI, comp3188minJ;
    Comparator comp3188(comp2650minVal, comp2650minI, comp2650minJ, comp2651minVal, comp2651minI, comp2651minJ, comp3188minVal, comp3188minI, comp3188minJ);
    wire [11:0] comp3189minVal;
    wire [5:0] comp3189minI, comp3189minJ;
    Comparator comp3189(comp2652minVal, comp2652minI, comp2652minJ, comp2653minVal, comp2653minI, comp2653minJ, comp3189minVal, comp3189minI, comp3189minJ);
    wire [11:0] comp3190minVal;
    wire [5:0] comp3190minI, comp3190minJ;
    Comparator comp3190(comp2654minVal, comp2654minI, comp2654minJ, comp2655minVal, comp2655minI, comp2655minJ, comp3190minVal, comp3190minI, comp3190minJ);
    wire [11:0] comp3191minVal;
    wire [5:0] comp3191minI, comp3191minJ;
    Comparator comp3191(comp2656minVal, comp2656minI, comp2656minJ, comp2657minVal, comp2657minI, comp2657minJ, comp3191minVal, comp3191minI, comp3191minJ);
    wire [11:0] comp3192minVal;
    wire [5:0] comp3192minI, comp3192minJ;
    Comparator comp3192(comp2658minVal, comp2658minI, comp2658minJ, comp2659minVal, comp2659minI, comp2659minJ, comp3192minVal, comp3192minI, comp3192minJ);
    wire [11:0] comp3193minVal;
    wire [5:0] comp3193minI, comp3193minJ;
    Comparator comp3193(comp2660minVal, comp2660minI, comp2660minJ, comp2661minVal, comp2661minI, comp2661minJ, comp3193minVal, comp3193minI, comp3193minJ);
    wire [11:0] comp3194minVal;
    wire [5:0] comp3194minI, comp3194minJ;
    Comparator comp3194(comp2662minVal, comp2662minI, comp2662minJ, comp2663minVal, comp2663minI, comp2663minJ, comp3194minVal, comp3194minI, comp3194minJ);
    wire [11:0] comp3195minVal;
    wire [5:0] comp3195minI, comp3195minJ;
    Comparator comp3195(comp2664minVal, comp2664minI, comp2664minJ, comp2665minVal, comp2665minI, comp2665minJ, comp3195minVal, comp3195minI, comp3195minJ);
    wire [11:0] comp3196minVal;
    wire [5:0] comp3196minI, comp3196minJ;
    Comparator comp3196(comp2666minVal, comp2666minI, comp2666minJ, comp2667minVal, comp2667minI, comp2667minJ, comp3196minVal, comp3196minI, comp3196minJ);
    wire [11:0] comp3197minVal;
    wire [5:0] comp3197minI, comp3197minJ;
    Comparator comp3197(comp2668minVal, comp2668minI, comp2668minJ, comp2669minVal, comp2669minI, comp2669minJ, comp3197minVal, comp3197minI, comp3197minJ);
    wire [11:0] comp3198minVal;
    wire [5:0] comp3198minI, comp3198minJ;
    Comparator comp3198(comp2670minVal, comp2670minI, comp2670minJ, comp2671minVal, comp2671minI, comp2671minJ, comp3198minVal, comp3198minI, comp3198minJ);
    wire [11:0] comp3199minVal;
    wire [5:0] comp3199minI, comp3199minJ;
    Comparator comp3199(comp2672minVal, comp2672minI, comp2672minJ, comp2673minVal, comp2673minI, comp2673minJ, comp3199minVal, comp3199minI, comp3199minJ);
    wire [11:0] comp3200minVal;
    wire [5:0] comp3200minI, comp3200minJ;
    Comparator comp3200(comp2674minVal, comp2674minI, comp2674minJ, comp2675minVal, comp2675minI, comp2675minJ, comp3200minVal, comp3200minI, comp3200minJ);
    wire [11:0] comp3201minVal;
    wire [5:0] comp3201minI, comp3201minJ;
    Comparator comp3201(comp2676minVal, comp2676minI, comp2676minJ, comp2677minVal, comp2677minI, comp2677minJ, comp3201minVal, comp3201minI, comp3201minJ);
    wire [11:0] comp3202minVal;
    wire [5:0] comp3202minI, comp3202minJ;
    Comparator comp3202(comp2678minVal, comp2678minI, comp2678minJ, comp2679minVal, comp2679minI, comp2679minJ, comp3202minVal, comp3202minI, comp3202minJ);
    wire [11:0] comp3203minVal;
    wire [5:0] comp3203minI, comp3203minJ;
    Comparator comp3203(comp2680minVal, comp2680minI, comp2680minJ, comp2681minVal, comp2681minI, comp2681minJ, comp3203minVal, comp3203minI, comp3203minJ);
    wire [11:0] comp3204minVal;
    wire [5:0] comp3204minI, comp3204minJ;
    Comparator comp3204(comp2682minVal, comp2682minI, comp2682minJ, comp2683minVal, comp2683minI, comp2683minJ, comp3204minVal, comp3204minI, comp3204minJ);
    wire [11:0] comp3205minVal;
    wire [5:0] comp3205minI, comp3205minJ;
    Comparator comp3205(comp2684minVal, comp2684minI, comp2684minJ, comp2685minVal, comp2685minI, comp2685minJ, comp3205minVal, comp3205minI, comp3205minJ);
    wire [11:0] comp3206minVal;
    wire [5:0] comp3206minI, comp3206minJ;
    Comparator comp3206(comp2686minVal, comp2686minI, comp2686minJ, comp2687minVal, comp2687minI, comp2687minJ, comp3206minVal, comp3206minI, comp3206minJ);
    wire [11:0] comp3207minVal;
    wire [5:0] comp3207minI, comp3207minJ;
    Comparator comp3207(comp2688minVal, comp2688minI, comp2688minJ, comp2689minVal, comp2689minI, comp2689minJ, comp3207minVal, comp3207minI, comp3207minJ);
    wire [11:0] comp3208minVal;
    wire [5:0] comp3208minI, comp3208minJ;
    Comparator comp3208(comp2690minVal, comp2690minI, comp2690minJ, comp2691minVal, comp2691minI, comp2691minJ, comp3208minVal, comp3208minI, comp3208minJ);
    wire [11:0] comp3209minVal;
    wire [5:0] comp3209minI, comp3209minJ;
    Comparator comp3209(comp2692minVal, comp2692minI, comp2692minJ, comp2693minVal, comp2693minI, comp2693minJ, comp3209minVal, comp3209minI, comp3209minJ);
    wire [11:0] comp3210minVal;
    wire [5:0] comp3210minI, comp3210minJ;
    Comparator comp3210(comp2694minVal, comp2694minI, comp2694minJ, comp2695minVal, comp2695minI, comp2695minJ, comp3210minVal, comp3210minI, comp3210minJ);
    wire [11:0] comp3211minVal;
    wire [5:0] comp3211minI, comp3211minJ;
    Comparator comp3211(comp2696minVal, comp2696minI, comp2696minJ, comp2697minVal, comp2697minI, comp2697minJ, comp3211minVal, comp3211minI, comp3211minJ);
    wire [11:0] comp3212minVal;
    wire [5:0] comp3212minI, comp3212minJ;
    Comparator comp3212(comp2698minVal, comp2698minI, comp2698minJ, comp2699minVal, comp2699minI, comp2699minJ, comp3212minVal, comp3212minI, comp3212minJ);
    wire [11:0] comp3213minVal;
    wire [5:0] comp3213minI, comp3213minJ;
    Comparator comp3213(comp2700minVal, comp2700minI, comp2700minJ, comp2701minVal, comp2701minI, comp2701minJ, comp3213minVal, comp3213minI, comp3213minJ);
    wire [11:0] comp3214minVal;
    wire [5:0] comp3214minI, comp3214minJ;
    Comparator comp3214(comp2702minVal, comp2702minI, comp2702minJ, comp2703minVal, comp2703minI, comp2703minJ, comp3214minVal, comp3214minI, comp3214minJ);
    wire [11:0] comp3215minVal;
    wire [5:0] comp3215minI, comp3215minJ;
    Comparator comp3215(comp2704minVal, comp2704minI, comp2704minJ, comp2705minVal, comp2705minI, comp2705minJ, comp3215minVal, comp3215minI, comp3215minJ);
    wire [11:0] comp3216minVal;
    wire [5:0] comp3216minI, comp3216minJ;
    Comparator comp3216(comp2706minVal, comp2706minI, comp2706minJ, comp2707minVal, comp2707minI, comp2707minJ, comp3216minVal, comp3216minI, comp3216minJ);
    wire [11:0] comp3217minVal;
    wire [5:0] comp3217minI, comp3217minJ;
    Comparator comp3217(comp2708minVal, comp2708minI, comp2708minJ, comp2709minVal, comp2709minI, comp2709minJ, comp3217minVal, comp3217minI, comp3217minJ);
    wire [11:0] comp3218minVal;
    wire [5:0] comp3218minI, comp3218minJ;
    Comparator comp3218(comp2710minVal, comp2710minI, comp2710minJ, comp2711minVal, comp2711minI, comp2711minJ, comp3218minVal, comp3218minI, comp3218minJ);
    wire [11:0] comp3219minVal;
    wire [5:0] comp3219minI, comp3219minJ;
    Comparator comp3219(comp2712minVal, comp2712minI, comp2712minJ, comp2713minVal, comp2713minI, comp2713minJ, comp3219minVal, comp3219minI, comp3219minJ);
    wire [11:0] comp3220minVal;
    wire [5:0] comp3220minI, comp3220minJ;
    Comparator comp3220(comp2714minVal, comp2714minI, comp2714minJ, comp2715minVal, comp2715minI, comp2715minJ, comp3220minVal, comp3220minI, comp3220minJ);
    wire [11:0] comp3221minVal;
    wire [5:0] comp3221minI, comp3221minJ;
    Comparator comp3221(comp2716minVal, comp2716minI, comp2716minJ, comp2717minVal, comp2717minI, comp2717minJ, comp3221minVal, comp3221minI, comp3221minJ);
    wire [11:0] comp3222minVal;
    wire [5:0] comp3222minI, comp3222minJ;
    Comparator comp3222(comp2718minVal, comp2718minI, comp2718minJ, comp2719minVal, comp2719minI, comp2719minJ, comp3222minVal, comp3222minI, comp3222minJ);
    wire [11:0] comp3223minVal;
    wire [5:0] comp3223minI, comp3223minJ;
    Comparator comp3223(comp2720minVal, comp2720minI, comp2720minJ, comp2721minVal, comp2721minI, comp2721minJ, comp3223minVal, comp3223minI, comp3223minJ);
    wire [11:0] comp3224minVal;
    wire [5:0] comp3224minI, comp3224minJ;
    Comparator comp3224(comp2722minVal, comp2722minI, comp2722minJ, comp2723minVal, comp2723minI, comp2723minJ, comp3224minVal, comp3224minI, comp3224minJ);
    wire [11:0] comp3225minVal;
    wire [5:0] comp3225minI, comp3225minJ;
    Comparator comp3225(comp2724minVal, comp2724minI, comp2724minJ, comp2725minVal, comp2725minI, comp2725minJ, comp3225minVal, comp3225minI, comp3225minJ);
    wire [11:0] comp3226minVal;
    wire [5:0] comp3226minI, comp3226minJ;
    Comparator comp3226(comp2726minVal, comp2726minI, comp2726minJ, comp2727minVal, comp2727minI, comp2727minJ, comp3226minVal, comp3226minI, comp3226minJ);
    wire [11:0] comp3227minVal;
    wire [5:0] comp3227minI, comp3227minJ;
    Comparator comp3227(comp2728minVal, comp2728minI, comp2728minJ, comp2729minVal, comp2729minI, comp2729minJ, comp3227minVal, comp3227minI, comp3227minJ);
    wire [11:0] comp3228minVal;
    wire [5:0] comp3228minI, comp3228minJ;
    Comparator comp3228(comp2730minVal, comp2730minI, comp2730minJ, comp2731minVal, comp2731minI, comp2731minJ, comp3228minVal, comp3228minI, comp3228minJ);
    wire [11:0] comp3229minVal;
    wire [5:0] comp3229minI, comp3229minJ;
    Comparator comp3229(comp2732minVal, comp2732minI, comp2732minJ, comp2733minVal, comp2733minI, comp2733minJ, comp3229minVal, comp3229minI, comp3229minJ);
    wire [11:0] comp3230minVal;
    wire [5:0] comp3230minI, comp3230minJ;
    Comparator comp3230(comp2734minVal, comp2734minI, comp2734minJ, comp2735minVal, comp2735minI, comp2735minJ, comp3230minVal, comp3230minI, comp3230minJ);
    wire [11:0] comp3231minVal;
    wire [5:0] comp3231minI, comp3231minJ;
    Comparator comp3231(comp2736minVal, comp2736minI, comp2736minJ, comp2737minVal, comp2737minI, comp2737minJ, comp3231minVal, comp3231minI, comp3231minJ);
    wire [11:0] comp3232minVal;
    wire [5:0] comp3232minI, comp3232minJ;
    Comparator comp3232(comp2738minVal, comp2738minI, comp2738minJ, comp2739minVal, comp2739minI, comp2739minJ, comp3232minVal, comp3232minI, comp3232minJ);
    wire [11:0] comp3233minVal;
    wire [5:0] comp3233minI, comp3233minJ;
    Comparator comp3233(comp2740minVal, comp2740minI, comp2740minJ, comp2741minVal, comp2741minI, comp2741minJ, comp3233minVal, comp3233minI, comp3233minJ);
    wire [11:0] comp3234minVal;
    wire [5:0] comp3234minI, comp3234minJ;
    Comparator comp3234(comp2742minVal, comp2742minI, comp2742minJ, comp2743minVal, comp2743minI, comp2743minJ, comp3234minVal, comp3234minI, comp3234minJ);
    wire [11:0] comp3235minVal;
    wire [5:0] comp3235minI, comp3235minJ;
    Comparator comp3235(comp2744minVal, comp2744minI, comp2744minJ, comp2745minVal, comp2745minI, comp2745minJ, comp3235minVal, comp3235minI, comp3235minJ);
    wire [11:0] comp3236minVal;
    wire [5:0] comp3236minI, comp3236minJ;
    Comparator comp3236(comp2746minVal, comp2746minI, comp2746minJ, comp2747minVal, comp2747minI, comp2747minJ, comp3236minVal, comp3236minI, comp3236minJ);
    wire [11:0] comp3237minVal;
    wire [5:0] comp3237minI, comp3237minJ;
    Comparator comp3237(comp2748minVal, comp2748minI, comp2748minJ, comp2749minVal, comp2749minI, comp2749minJ, comp3237minVal, comp3237minI, comp3237minJ);
    wire [11:0] comp3238minVal;
    wire [5:0] comp3238minI, comp3238minJ;
    Comparator comp3238(comp2750minVal, comp2750minI, comp2750minJ, comp2751minVal, comp2751minI, comp2751minJ, comp3238minVal, comp3238minI, comp3238minJ);
    wire [11:0] comp3239minVal;
    wire [5:0] comp3239minI, comp3239minJ;
    Comparator comp3239(comp2752minVal, comp2752minI, comp2752minJ, comp2753minVal, comp2753minI, comp2753minJ, comp3239minVal, comp3239minI, comp3239minJ);
    wire [11:0] comp3240minVal;
    wire [5:0] comp3240minI, comp3240minJ;
    Comparator comp3240(comp2754minVal, comp2754minI, comp2754minJ, comp2755minVal, comp2755minI, comp2755minJ, comp3240minVal, comp3240minI, comp3240minJ);
    wire [11:0] comp3241minVal;
    wire [5:0] comp3241minI, comp3241minJ;
    Comparator comp3241(comp2756minVal, comp2756minI, comp2756minJ, comp2757minVal, comp2757minI, comp2757minJ, comp3241minVal, comp3241minI, comp3241minJ);
    wire [11:0] comp3242minVal;
    wire [5:0] comp3242minI, comp3242minJ;
    Comparator comp3242(comp2758minVal, comp2758minI, comp2758minJ, comp2759minVal, comp2759minI, comp2759minJ, comp3242minVal, comp3242minI, comp3242minJ);
    wire [11:0] comp3243minVal;
    wire [5:0] comp3243minI, comp3243minJ;
    Comparator comp3243(comp2760minVal, comp2760minI, comp2760minJ, comp2761minVal, comp2761minI, comp2761minJ, comp3243minVal, comp3243minI, comp3243minJ);
    wire [11:0] comp3244minVal;
    wire [5:0] comp3244minI, comp3244minJ;
    Comparator comp3244(comp2762minVal, comp2762minI, comp2762minJ, comp2763minVal, comp2763minI, comp2763minJ, comp3244minVal, comp3244minI, comp3244minJ);
    wire [11:0] comp3245minVal;
    wire [5:0] comp3245minI, comp3245minJ;
    Comparator comp3245(comp2764minVal, comp2764minI, comp2764minJ, comp2765minVal, comp2765minI, comp2765minJ, comp3245minVal, comp3245minI, comp3245minJ);
    wire [11:0] comp3246minVal;
    wire [5:0] comp3246minI, comp3246minJ;
    Comparator comp3246(comp2766minVal, comp2766minI, comp2766minJ, comp2767minVal, comp2767minI, comp2767minJ, comp3246minVal, comp3246minI, comp3246minJ);
    wire [11:0] comp3247minVal;
    wire [5:0] comp3247minI, comp3247minJ;
    Comparator comp3247(comp2768minVal, comp2768minI, comp2768minJ, comp2769minVal, comp2769minI, comp2769minJ, comp3247minVal, comp3247minI, comp3247minJ);
    wire [11:0] comp3248minVal;
    wire [5:0] comp3248minI, comp3248minJ;
    Comparator comp3248(comp2770minVal, comp2770minI, comp2770minJ, comp2771minVal, comp2771minI, comp2771minJ, comp3248minVal, comp3248minI, comp3248minJ);
    wire [11:0] comp3249minVal;
    wire [5:0] comp3249minI, comp3249minJ;
    Comparator comp3249(comp2772minVal, comp2772minI, comp2772minJ, comp2773minVal, comp2773minI, comp2773minJ, comp3249minVal, comp3249minI, comp3249minJ);
    wire [11:0] comp3250minVal;
    wire [5:0] comp3250minI, comp3250minJ;
    Comparator comp3250(comp2774minVal, comp2774minI, comp2774minJ, comp2775minVal, comp2775minI, comp2775minJ, comp3250minVal, comp3250minI, comp3250minJ);
    wire [11:0] comp3251minVal;
    wire [5:0] comp3251minI, comp3251minJ;
    Comparator comp3251(comp2776minVal, comp2776minI, comp2776minJ, comp2777minVal, comp2777minI, comp2777minJ, comp3251minVal, comp3251minI, comp3251minJ);
    wire [11:0] comp3252minVal;
    wire [5:0] comp3252minI, comp3252minJ;
    Comparator comp3252(comp2778minVal, comp2778minI, comp2778minJ, comp2779minVal, comp2779minI, comp2779minJ, comp3252minVal, comp3252minI, comp3252minJ);
    wire [11:0] comp3253minVal;
    wire [5:0] comp3253minI, comp3253minJ;
    Comparator comp3253(comp2780minVal, comp2780minI, comp2780minJ, comp2781minVal, comp2781minI, comp2781minJ, comp3253minVal, comp3253minI, comp3253minJ);
    wire [11:0] comp3254minVal;
    wire [5:0] comp3254minI, comp3254minJ;
    Comparator comp3254(comp2782minVal, comp2782minI, comp2782minJ, comp2783minVal, comp2783minI, comp2783minJ, comp3254minVal, comp3254minI, comp3254minJ);
    wire [11:0] comp3255minVal;
    wire [5:0] comp3255minI, comp3255minJ;
    Comparator comp3255(comp2784minVal, comp2784minI, comp2784minJ, comp2785minVal, comp2785minI, comp2785minJ, comp3255minVal, comp3255minI, comp3255minJ);
    wire [11:0] comp3256minVal;
    wire [5:0] comp3256minI, comp3256minJ;
    Comparator comp3256(comp2786minVal, comp2786minI, comp2786minJ, comp2787minVal, comp2787minI, comp2787minJ, comp3256minVal, comp3256minI, comp3256minJ);
    wire [11:0] comp3257minVal;
    wire [5:0] comp3257minI, comp3257minJ;
    Comparator comp3257(comp2788minVal, comp2788minI, comp2788minJ, comp2789minVal, comp2789minI, comp2789minJ, comp3257minVal, comp3257minI, comp3257minJ);
    wire [11:0] comp3258minVal;
    wire [5:0] comp3258minI, comp3258minJ;
    Comparator comp3258(comp2790minVal, comp2790minI, comp2790minJ, comp2791minVal, comp2791minI, comp2791minJ, comp3258minVal, comp3258minI, comp3258minJ);
    wire [11:0] comp3259minVal;
    wire [5:0] comp3259minI, comp3259minJ;
    Comparator comp3259(comp2792minVal, comp2792minI, comp2792minJ, comp2793minVal, comp2793minI, comp2793minJ, comp3259minVal, comp3259minI, comp3259minJ);
    wire [11:0] comp3260minVal;
    wire [5:0] comp3260minI, comp3260minJ;
    Comparator comp3260(comp2794minVal, comp2794minI, comp2794minJ, comp2795minVal, comp2795minI, comp2795minJ, comp3260minVal, comp3260minI, comp3260minJ);
    wire [11:0] comp3261minVal;
    wire [5:0] comp3261minI, comp3261minJ;
    Comparator comp3261(comp2796minVal, comp2796minI, comp2796minJ, comp2797minVal, comp2797minI, comp2797minJ, comp3261minVal, comp3261minI, comp3261minJ);
    wire [11:0] comp3262minVal;
    wire [5:0] comp3262minI, comp3262minJ;
    Comparator comp3262(comp2798minVal, comp2798minI, comp2798minJ, comp2799minVal, comp2799minI, comp2799minJ, comp3262minVal, comp3262minI, comp3262minJ);
    wire [11:0] comp3263minVal;
    wire [5:0] comp3263minI, comp3263minJ;
    Comparator comp3263(comp2800minVal, comp2800minI, comp2800minJ, comp2801minVal, comp2801minI, comp2801minJ, comp3263minVal, comp3263minI, comp3263minJ);
    wire [11:0] comp3264minVal;
    wire [5:0] comp3264minI, comp3264minJ;
    Comparator comp3264(comp2802minVal, comp2802minI, comp2802minJ, comp2803minVal, comp2803minI, comp2803minJ, comp3264minVal, comp3264minI, comp3264minJ);
    wire [11:0] comp3265minVal;
    wire [5:0] comp3265minI, comp3265minJ;
    Comparator comp3265(comp2804minVal, comp2804minI, comp2804minJ, comp2805minVal, comp2805minI, comp2805minJ, comp3265minVal, comp3265minI, comp3265minJ);
    wire [11:0] comp3266minVal;
    wire [5:0] comp3266minI, comp3266minJ;
    Comparator comp3266(comp2806minVal, comp2806minI, comp2806minJ, comp2807minVal, comp2807minI, comp2807minJ, comp3266minVal, comp3266minI, comp3266minJ);
    wire [11:0] comp3267minVal;
    wire [5:0] comp3267minI, comp3267minJ;
    Comparator comp3267(comp2808minVal, comp2808minI, comp2808minJ, comp2809minVal, comp2809minI, comp2809minJ, comp3267minVal, comp3267minI, comp3267minJ);
    wire [11:0] comp3268minVal;
    wire [5:0] comp3268minI, comp3268minJ;
    Comparator comp3268(comp2810minVal, comp2810minI, comp2810minJ, comp2811minVal, comp2811minI, comp2811minJ, comp3268minVal, comp3268minI, comp3268minJ);
    wire [11:0] comp3269minVal;
    wire [5:0] comp3269minI, comp3269minJ;
    Comparator comp3269(comp2812minVal, comp2812minI, comp2812minJ, comp2813minVal, comp2813minI, comp2813minJ, comp3269minVal, comp3269minI, comp3269minJ);
    wire [11:0] comp3270minVal;
    wire [5:0] comp3270minI, comp3270minJ;
    Comparator comp3270(comp2814minVal, comp2814minI, comp2814minJ, comp2815minVal, comp2815minI, comp2815minJ, comp3270minVal, comp3270minI, comp3270minJ);
    wire [11:0] comp3271minVal;
    wire [5:0] comp3271minI, comp3271minJ;
    Comparator comp3271(comp2816minVal, comp2816minI, comp2816minJ, comp2817minVal, comp2817minI, comp2817minJ, comp3271minVal, comp3271minI, comp3271minJ);
    wire [11:0] comp3272minVal;
    wire [5:0] comp3272minI, comp3272minJ;
    Comparator comp3272(comp2818minVal, comp2818minI, comp2818minJ, comp2819minVal, comp2819minI, comp2819minJ, comp3272minVal, comp3272minI, comp3272minJ);
    wire [11:0] comp3273minVal;
    wire [5:0] comp3273minI, comp3273minJ;
    Comparator comp3273(comp2820minVal, comp2820minI, comp2820minJ, comp2821minVal, comp2821minI, comp2821minJ, comp3273minVal, comp3273minI, comp3273minJ);
    wire [11:0] comp3274minVal;
    wire [5:0] comp3274minI, comp3274minJ;
    Comparator comp3274(comp2822minVal, comp2822minI, comp2822minJ, comp2823minVal, comp2823minI, comp2823minJ, comp3274minVal, comp3274minI, comp3274minJ);
    wire [11:0] comp3275minVal;
    wire [5:0] comp3275minI, comp3275minJ;
    Comparator comp3275(comp2824minVal, comp2824minI, comp2824minJ, comp2825minVal, comp2825minI, comp2825minJ, comp3275minVal, comp3275minI, comp3275minJ);
    wire [11:0] comp3276minVal;
    wire [5:0] comp3276minI, comp3276minJ;
    Comparator comp3276(comp2826minVal, comp2826minI, comp2826minJ, comp2827minVal, comp2827minI, comp2827minJ, comp3276minVal, comp3276minI, comp3276minJ);
    wire [11:0] comp3277minVal;
    wire [5:0] comp3277minI, comp3277minJ;
    Comparator comp3277(comp2828minVal, comp2828minI, comp2828minJ, comp2829minVal, comp2829minI, comp2829minJ, comp3277minVal, comp3277minI, comp3277minJ);
    wire [11:0] comp3278minVal;
    wire [5:0] comp3278minI, comp3278minJ;
    Comparator comp3278(comp2830minVal, comp2830minI, comp2830minJ, comp2831minVal, comp2831minI, comp2831minJ, comp3278minVal, comp3278minI, comp3278minJ);
    wire [11:0] comp3279minVal;
    wire [5:0] comp3279minI, comp3279minJ;
    Comparator comp3279(comp2832minVal, comp2832minI, comp2832minJ, comp2833minVal, comp2833minI, comp2833minJ, comp3279minVal, comp3279minI, comp3279minJ);
    wire [11:0] comp3280minVal;
    wire [5:0] comp3280minI, comp3280minJ;
    Comparator comp3280(comp2834minVal, comp2834minI, comp2834minJ, comp2835minVal, comp2835minI, comp2835minJ, comp3280minVal, comp3280minI, comp3280minJ);
    wire [11:0] comp3281minVal;
    wire [5:0] comp3281minI, comp3281minJ;
    Comparator comp3281(comp2836minVal, comp2836minI, comp2836minJ, comp2837minVal, comp2837minI, comp2837minJ, comp3281minVal, comp3281minI, comp3281minJ);
    wire [11:0] comp3282minVal;
    wire [5:0] comp3282minI, comp3282minJ;
    Comparator comp3282(comp2838minVal, comp2838minI, comp2838minJ, comp2839minVal, comp2839minI, comp2839minJ, comp3282minVal, comp3282minI, comp3282minJ);
    wire [11:0] comp3283minVal;
    wire [5:0] comp3283minI, comp3283minJ;
    Comparator comp3283(comp2840minVal, comp2840minI, comp2840minJ, comp2841minVal, comp2841minI, comp2841minJ, comp3283minVal, comp3283minI, comp3283minJ);
    wire [11:0] comp3284minVal;
    wire [5:0] comp3284minI, comp3284minJ;
    Comparator comp3284(comp2842minVal, comp2842minI, comp2842minJ, comp2843minVal, comp2843minI, comp2843minJ, comp3284minVal, comp3284minI, comp3284minJ);
    wire [11:0] comp3285minVal;
    wire [5:0] comp3285minI, comp3285minJ;
    Comparator comp3285(comp2844minVal, comp2844minI, comp2844minJ, comp2845minVal, comp2845minI, comp2845minJ, comp3285minVal, comp3285minI, comp3285minJ);
    wire [11:0] comp3286minVal;
    wire [5:0] comp3286minI, comp3286minJ;
    Comparator comp3286(comp2846minVal, comp2846minI, comp2846minJ, comp2847minVal, comp2847minI, comp2847minJ, comp3286minVal, comp3286minI, comp3286minJ);
    wire [11:0] comp3287minVal;
    wire [5:0] comp3287minI, comp3287minJ;
    Comparator comp3287(comp2848minVal, comp2848minI, comp2848minJ, comp2849minVal, comp2849minI, comp2849minJ, comp3287minVal, comp3287minI, comp3287minJ);
    wire [11:0] comp3288minVal;
    wire [5:0] comp3288minI, comp3288minJ;
    Comparator comp3288(comp2850minVal, comp2850minI, comp2850minJ, comp2851minVal, comp2851minI, comp2851minJ, comp3288minVal, comp3288minI, comp3288minJ);
    wire [11:0] comp3289minVal;
    wire [5:0] comp3289minI, comp3289minJ;
    Comparator comp3289(comp2852minVal, comp2852minI, comp2852minJ, comp2853minVal, comp2853minI, comp2853minJ, comp3289minVal, comp3289minI, comp3289minJ);
    wire [11:0] comp3290minVal;
    wire [5:0] comp3290minI, comp3290minJ;
    Comparator comp3290(comp2854minVal, comp2854minI, comp2854minJ, comp2855minVal, comp2855minI, comp2855minJ, comp3290minVal, comp3290minI, comp3290minJ);
    wire [11:0] comp3291minVal;
    wire [5:0] comp3291minI, comp3291minJ;
    Comparator comp3291(comp2856minVal, comp2856minI, comp2856minJ, comp2857minVal, comp2857minI, comp2857minJ, comp3291minVal, comp3291minI, comp3291minJ);
    wire [11:0] comp3292minVal;
    wire [5:0] comp3292minI, comp3292minJ;
    Comparator comp3292(comp2858minVal, comp2858minI, comp2858minJ, comp2859minVal, comp2859minI, comp2859minJ, comp3292minVal, comp3292minI, comp3292minJ);
    wire [11:0] comp3293minVal;
    wire [5:0] comp3293minI, comp3293minJ;
    Comparator comp3293(comp2860minVal, comp2860minI, comp2860minJ, comp2861minVal, comp2861minI, comp2861minJ, comp3293minVal, comp3293minI, comp3293minJ);
    wire [11:0] comp3294minVal;
    wire [5:0] comp3294minI, comp3294minJ;
    Comparator comp3294(comp2862minVal, comp2862minI, comp2862minJ, comp2863minVal, comp2863minI, comp2863minJ, comp3294minVal, comp3294minI, comp3294minJ);
    wire [11:0] comp3295minVal;
    wire [5:0] comp3295minI, comp3295minJ;
    Comparator comp3295(comp2864minVal, comp2864minI, comp2864minJ, comp2865minVal, comp2865minI, comp2865minJ, comp3295minVal, comp3295minI, comp3295minJ);
    wire [11:0] comp3296minVal;
    wire [5:0] comp3296minI, comp3296minJ;
    Comparator comp3296(comp2866minVal, comp2866minI, comp2866minJ, comp2867minVal, comp2867minI, comp2867minJ, comp3296minVal, comp3296minI, comp3296minJ);
    wire [11:0] comp3297minVal;
    wire [5:0] comp3297minI, comp3297minJ;
    Comparator comp3297(comp2868minVal, comp2868minI, comp2868minJ, comp2869minVal, comp2869minI, comp2869minJ, comp3297minVal, comp3297minI, comp3297minJ);
    wire [11:0] comp3298minVal;
    wire [5:0] comp3298minI, comp3298minJ;
    Comparator comp3298(comp2870minVal, comp2870minI, comp2870minJ, comp2871minVal, comp2871minI, comp2871minJ, comp3298minVal, comp3298minI, comp3298minJ);
    wire [11:0] comp3299minVal;
    wire [5:0] comp3299minI, comp3299minJ;
    Comparator comp3299(comp2872minVal, comp2872minI, comp2872minJ, comp2873minVal, comp2873minI, comp2873minJ, comp3299minVal, comp3299minI, comp3299minJ);
    wire [11:0] comp3300minVal;
    wire [5:0] comp3300minI, comp3300minJ;
    Comparator comp3300(comp2874minVal, comp2874minI, comp2874minJ, comp2875minVal, comp2875minI, comp2875minJ, comp3300minVal, comp3300minI, comp3300minJ);
    wire [11:0] comp3301minVal;
    wire [5:0] comp3301minI, comp3301minJ;
    Comparator comp3301(comp2876minVal, comp2876minI, comp2876minJ, comp2877minVal, comp2877minI, comp2877minJ, comp3301minVal, comp3301minI, comp3301minJ);
    wire [11:0] comp3302minVal;
    wire [5:0] comp3302minI, comp3302minJ;
    Comparator comp3302(comp2878minVal, comp2878minI, comp2878minJ, comp2879minVal, comp2879minI, comp2879minJ, comp3302minVal, comp3302minI, comp3302minJ);
    wire [11:0] comp3303minVal;
    wire [5:0] comp3303minI, comp3303minJ;
    Comparator comp3303(comp2880minVal, comp2880minI, comp2880minJ, comp2881minVal, comp2881minI, comp2881minJ, comp3303minVal, comp3303minI, comp3303minJ);
    wire [11:0] comp3304minVal;
    wire [5:0] comp3304minI, comp3304minJ;
    Comparator comp3304(comp2882minVal, comp2882minI, comp2882minJ, comp2883minVal, comp2883minI, comp2883minJ, comp3304minVal, comp3304minI, comp3304minJ);
    wire [11:0] comp3305minVal;
    wire [5:0] comp3305minI, comp3305minJ;
    Comparator comp3305(comp2884minVal, comp2884minI, comp2884minJ, comp2885minVal, comp2885minI, comp2885minJ, comp3305minVal, comp3305minI, comp3305minJ);
    wire [11:0] comp3306minVal;
    wire [5:0] comp3306minI, comp3306minJ;
    Comparator comp3306(comp2886minVal, comp2886minI, comp2886minJ, comp2887minVal, comp2887minI, comp2887minJ, comp3306minVal, comp3306minI, comp3306minJ);
    wire [11:0] comp3307minVal;
    wire [5:0] comp3307minI, comp3307minJ;
    Comparator comp3307(comp2888minVal, comp2888minI, comp2888minJ, comp2889minVal, comp2889minI, comp2889minJ, comp3307minVal, comp3307minI, comp3307minJ);
    wire [11:0] comp3308minVal;
    wire [5:0] comp3308minI, comp3308minJ;
    Comparator comp3308(comp2890minVal, comp2890minI, comp2890minJ, comp2891minVal, comp2891minI, comp2891minJ, comp3308minVal, comp3308minI, comp3308minJ);
    wire [11:0] comp3309minVal;
    wire [5:0] comp3309minI, comp3309minJ;
    Comparator comp3309(comp2892minVal, comp2892minI, comp2892minJ, comp2893minVal, comp2893minI, comp2893minJ, comp3309minVal, comp3309minI, comp3309minJ);
    wire [11:0] comp3310minVal;
    wire [5:0] comp3310minI, comp3310minJ;
    Comparator comp3310(comp2894minVal, comp2894minI, comp2894minJ, comp2895minVal, comp2895minI, comp2895minJ, comp3310minVal, comp3310minI, comp3310minJ);
    wire [11:0] comp3311minVal;
    wire [5:0] comp3311minI, comp3311minJ;
    Comparator comp3311(comp2896minVal, comp2896minI, comp2896minJ, comp2897minVal, comp2897minI, comp2897minJ, comp3311minVal, comp3311minI, comp3311minJ);
    wire [11:0] comp3312minVal;
    wire [5:0] comp3312minI, comp3312minJ;
    Comparator comp3312(comp2898minVal, comp2898minI, comp2898minJ, comp2899minVal, comp2899minI, comp2899minJ, comp3312minVal, comp3312minI, comp3312minJ);
    wire [11:0] comp3313minVal;
    wire [5:0] comp3313minI, comp3313minJ;
    Comparator comp3313(comp2900minVal, comp2900minI, comp2900minJ, comp2901minVal, comp2901minI, comp2901minJ, comp3313minVal, comp3313minI, comp3313minJ);
    wire [11:0] comp3314minVal;
    wire [5:0] comp3314minI, comp3314minJ;
    Comparator comp3314(comp2902minVal, comp2902minI, comp2902minJ, comp2903minVal, comp2903minI, comp2903minJ, comp3314minVal, comp3314minI, comp3314minJ);
    wire [11:0] comp3315minVal;
    wire [5:0] comp3315minI, comp3315minJ;
    Comparator comp3315(comp2904minVal, comp2904minI, comp2904minJ, comp2905minVal, comp2905minI, comp2905minJ, comp3315minVal, comp3315minI, comp3315minJ);
    wire [11:0] comp3316minVal;
    wire [5:0] comp3316minI, comp3316minJ;
    Comparator comp3316(comp2906minVal, comp2906minI, comp2906minJ, comp2907minVal, comp2907minI, comp2907minJ, comp3316minVal, comp3316minI, comp3316minJ);
    wire [11:0] comp3317minVal;
    wire [5:0] comp3317minI, comp3317minJ;
    Comparator comp3317(comp2908minVal, comp2908minI, comp2908minJ, comp2909minVal, comp2909minI, comp2909minJ, comp3317minVal, comp3317minI, comp3317minJ);
    wire [11:0] comp3318minVal;
    wire [5:0] comp3318minI, comp3318minJ;
    Comparator comp3318(comp2910minVal, comp2910minI, comp2910minJ, comp2911minVal, comp2911minI, comp2911minJ, comp3318minVal, comp3318minI, comp3318minJ);
    wire [11:0] comp3319minVal;
    wire [5:0] comp3319minI, comp3319minJ;
    Comparator comp3319(comp2912minVal, comp2912minI, comp2912minJ, comp2913minVal, comp2913minI, comp2913minJ, comp3319minVal, comp3319minI, comp3319minJ);
    wire [11:0] comp3320minVal;
    wire [5:0] comp3320minI, comp3320minJ;
    Comparator comp3320(comp2914minVal, comp2914minI, comp2914minJ, comp2915minVal, comp2915minI, comp2915minJ, comp3320minVal, comp3320minI, comp3320minJ);
    wire [11:0] comp3321minVal;
    wire [5:0] comp3321minI, comp3321minJ;
    Comparator comp3321(comp2916minVal, comp2916minI, comp2916minJ, comp2917minVal, comp2917minI, comp2917minJ, comp3321minVal, comp3321minI, comp3321minJ);
    wire [11:0] comp3322minVal;
    wire [5:0] comp3322minI, comp3322minJ;
    Comparator comp3322(comp2918minVal, comp2918minI, comp2918minJ, comp2919minVal, comp2919minI, comp2919minJ, comp3322minVal, comp3322minI, comp3322minJ);
    wire [11:0] comp3323minVal;
    wire [5:0] comp3323minI, comp3323minJ;
    Comparator comp3323(comp2920minVal, comp2920minI, comp2920minJ, comp2921minVal, comp2921minI, comp2921minJ, comp3323minVal, comp3323minI, comp3323minJ);
    wire [11:0] comp3324minVal;
    wire [5:0] comp3324minI, comp3324minJ;
    Comparator comp3324(comp2922minVal, comp2922minI, comp2922minJ, comp2923minVal, comp2923minI, comp2923minJ, comp3324minVal, comp3324minI, comp3324minJ);
    wire [11:0] comp3325minVal;
    wire [5:0] comp3325minI, comp3325minJ;
    Comparator comp3325(comp2924minVal, comp2924minI, comp2924minJ, comp2925minVal, comp2925minI, comp2925minJ, comp3325minVal, comp3325minI, comp3325minJ);
    wire [11:0] comp3326minVal;
    wire [5:0] comp3326minI, comp3326minJ;
    Comparator comp3326(comp2926minVal, comp2926minI, comp2926minJ, comp2927minVal, comp2927minI, comp2927minJ, comp3326minVal, comp3326minI, comp3326minJ);
    wire [11:0] comp3327minVal;
    wire [5:0] comp3327minI, comp3327minJ;
    Comparator comp3327(comp2928minVal, comp2928minI, comp2928minJ, comp2929minVal, comp2929minI, comp2929minJ, comp3327minVal, comp3327minI, comp3327minJ);
    wire [11:0] comp3328minVal;
    wire [5:0] comp3328minI, comp3328minJ;
    Comparator comp3328(comp2930minVal, comp2930minI, comp2930minJ, comp2931minVal, comp2931minI, comp2931minJ, comp3328minVal, comp3328minI, comp3328minJ);
    wire [11:0] comp3329minVal;
    wire [5:0] comp3329minI, comp3329minJ;
    Comparator comp3329(comp2932minVal, comp2932minI, comp2932minJ, comp2933minVal, comp2933minI, comp2933minJ, comp3329minVal, comp3329minI, comp3329minJ);
    wire [11:0] comp3330minVal;
    wire [5:0] comp3330minI, comp3330minJ;
    Comparator comp3330(comp2934minVal, comp2934minI, comp2934minJ, comp2935minVal, comp2935minI, comp2935minJ, comp3330minVal, comp3330minI, comp3330minJ);
    wire [11:0] comp3331minVal;
    wire [5:0] comp3331minI, comp3331minJ;
    Comparator comp3331(comp2936minVal, comp2936minI, comp2936minJ, comp2937minVal, comp2937minI, comp2937minJ, comp3331minVal, comp3331minI, comp3331minJ);
    wire [11:0] comp3332minVal;
    wire [5:0] comp3332minI, comp3332minJ;
    Comparator comp3332(comp2938minVal, comp2938minI, comp2938minJ, comp2939minVal, comp2939minI, comp2939minJ, comp3332minVal, comp3332minI, comp3332minJ);
    wire [11:0] comp3333minVal;
    wire [5:0] comp3333minI, comp3333minJ;
    Comparator comp3333(comp2940minVal, comp2940minI, comp2940minJ, comp2941minVal, comp2941minI, comp2941minJ, comp3333minVal, comp3333minI, comp3333minJ);
    wire [11:0] comp3334minVal;
    wire [5:0] comp3334minI, comp3334minJ;
    Comparator comp3334(comp2942minVal, comp2942minI, comp2942minJ, comp2943minVal, comp2943minI, comp2943minJ, comp3334minVal, comp3334minI, comp3334minJ);
    wire [11:0] comp3335minVal;
    wire [5:0] comp3335minI, comp3335minJ;
    Comparator comp3335(comp2944minVal, comp2944minI, comp2944minJ, comp2945minVal, comp2945minI, comp2945minJ, comp3335minVal, comp3335minI, comp3335minJ);
    wire [11:0] comp3336minVal;
    wire [5:0] comp3336minI, comp3336minJ;
    Comparator comp3336(comp2946minVal, comp2946minI, comp2946minJ, comp2947minVal, comp2947minI, comp2947minJ, comp3336minVal, comp3336minI, comp3336minJ);
    wire [11:0] comp3337minVal;
    wire [5:0] comp3337minI, comp3337minJ;
    Comparator comp3337(comp2948minVal, comp2948minI, comp2948minJ, comp2949minVal, comp2949minI, comp2949minJ, comp3337minVal, comp3337minI, comp3337minJ);
    wire [11:0] comp3338minVal;
    wire [5:0] comp3338minI, comp3338minJ;
    Comparator comp3338(comp2950minVal, comp2950minI, comp2950minJ, comp2951minVal, comp2951minI, comp2951minJ, comp3338minVal, comp3338minI, comp3338minJ);
    wire [11:0] comp3339minVal;
    wire [5:0] comp3339minI, comp3339minJ;
    Comparator comp3339(comp2952minVal, comp2952minI, comp2952minJ, comp2953minVal, comp2953minI, comp2953minJ, comp3339minVal, comp3339minI, comp3339minJ);
    wire [11:0] comp3340minVal;
    wire [5:0] comp3340minI, comp3340minJ;
    Comparator comp3340(comp2954minVal, comp2954minI, comp2954minJ, comp2955minVal, comp2955minI, comp2955minJ, comp3340minVal, comp3340minI, comp3340minJ);
    wire [11:0] comp3341minVal;
    wire [5:0] comp3341minI, comp3341minJ;
    Comparator comp3341(comp2956minVal, comp2956minI, comp2956minJ, comp2957minVal, comp2957minI, comp2957minJ, comp3341minVal, comp3341minI, comp3341minJ);
    wire [11:0] comp3342minVal;
    wire [5:0] comp3342minI, comp3342minJ;
    Comparator comp3342(comp2958minVal, comp2958minI, comp2958minJ, comp2959minVal, comp2959minI, comp2959minJ, comp3342minVal, comp3342minI, comp3342minJ);
    wire [11:0] comp3343minVal;
    wire [5:0] comp3343minI, comp3343minJ;
    Comparator comp3343(comp2960minVal, comp2960minI, comp2960minJ, comp2961minVal, comp2961minI, comp2961minJ, comp3343minVal, comp3343minI, comp3343minJ);
    wire [11:0] comp3344minVal;
    wire [5:0] comp3344minI, comp3344minJ;
    Comparator comp3344(comp2962minVal, comp2962minI, comp2962minJ, comp2963minVal, comp2963minI, comp2963minJ, comp3344minVal, comp3344minI, comp3344minJ);
    wire [11:0] comp3345minVal;
    wire [5:0] comp3345minI, comp3345minJ;
    Comparator comp3345(comp2964minVal, comp2964minI, comp2964minJ, comp2965minVal, comp2965minI, comp2965minJ, comp3345minVal, comp3345minI, comp3345minJ);
    wire [11:0] comp3346minVal;
    wire [5:0] comp3346minI, comp3346minJ;
    Comparator comp3346(comp2966minVal, comp2966minI, comp2966minJ, comp2967minVal, comp2967minI, comp2967minJ, comp3346minVal, comp3346minI, comp3346minJ);
    wire [11:0] comp3347minVal;
    wire [5:0] comp3347minI, comp3347minJ;
    Comparator comp3347(comp2968minVal, comp2968minI, comp2968minJ, comp2969minVal, comp2969minI, comp2969minJ, comp3347minVal, comp3347minI, comp3347minJ);
    wire [11:0] comp3348minVal;
    wire [5:0] comp3348minI, comp3348minJ;
    Comparator comp3348(comp2970minVal, comp2970minI, comp2970minJ, comp2971minVal, comp2971minI, comp2971minJ, comp3348minVal, comp3348minI, comp3348minJ);
    wire [11:0] comp3349minVal;
    wire [5:0] comp3349minI, comp3349minJ;
    Comparator comp3349(comp2972minVal, comp2972minI, comp2972minJ, comp2973minVal, comp2973minI, comp2973minJ, comp3349minVal, comp3349minI, comp3349minJ);
    wire [11:0] comp3350minVal;
    wire [5:0] comp3350minI, comp3350minJ;
    Comparator comp3350(comp2974minVal, comp2974minI, comp2974minJ, comp2975minVal, comp2975minI, comp2975minJ, comp3350minVal, comp3350minI, comp3350minJ);
    wire [11:0] comp3351minVal;
    wire [5:0] comp3351minI, comp3351minJ;
    Comparator comp3351(comp2976minVal, comp2976minI, comp2976minJ, comp2977minVal, comp2977minI, comp2977minJ, comp3351minVal, comp3351minI, comp3351minJ);
    wire [11:0] comp3352minVal;
    wire [5:0] comp3352minI, comp3352minJ;
    Comparator comp3352(comp2978minVal, comp2978minI, comp2978minJ, comp2979minVal, comp2979minI, comp2979minJ, comp3352minVal, comp3352minI, comp3352minJ);
    wire [11:0] comp3353minVal;
    wire [5:0] comp3353minI, comp3353minJ;
    Comparator comp3353(comp2980minVal, comp2980minI, comp2980minJ, comp2981minVal, comp2981minI, comp2981minJ, comp3353minVal, comp3353minI, comp3353minJ);
    wire [11:0] comp3354minVal;
    wire [5:0] comp3354minI, comp3354minJ;
    Comparator comp3354(comp2982minVal, comp2982minI, comp2982minJ, comp2983minVal, comp2983minI, comp2983minJ, comp3354minVal, comp3354minI, comp3354minJ);
    wire [11:0] comp3355minVal;
    wire [5:0] comp3355minI, comp3355minJ;
    Comparator comp3355(comp2984minVal, comp2984minI, comp2984minJ, comp2985minVal, comp2985minI, comp2985minJ, comp3355minVal, comp3355minI, comp3355minJ);
    wire [11:0] comp3356minVal;
    wire [5:0] comp3356minI, comp3356minJ;
    Comparator comp3356(comp2986minVal, comp2986minI, comp2986minJ, comp2987minVal, comp2987minI, comp2987minJ, comp3356minVal, comp3356minI, comp3356minJ);
    wire [11:0] comp3357minVal;
    wire [5:0] comp3357minI, comp3357minJ;
    Comparator comp3357(comp2988minVal, comp2988minI, comp2988minJ, comp2989minVal, comp2989minI, comp2989minJ, comp3357minVal, comp3357minI, comp3357minJ);
    wire [11:0] comp3358minVal;
    wire [5:0] comp3358minI, comp3358minJ;
    Comparator comp3358(comp2990minVal, comp2990minI, comp2990minJ, comp2991minVal, comp2991minI, comp2991minJ, comp3358minVal, comp3358minI, comp3358minJ);
    wire [11:0] comp3359minVal;
    wire [5:0] comp3359minI, comp3359minJ;
    Comparator comp3359(comp2992minVal, comp2992minI, comp2992minJ, comp2993minVal, comp2993minI, comp2993minJ, comp3359minVal, comp3359minI, comp3359minJ);
    wire [11:0] comp3360minVal;
    wire [5:0] comp3360minI, comp3360minJ;
    Comparator comp3360(comp2994minVal, comp2994minI, comp2994minJ, comp2995minVal, comp2995minI, comp2995minJ, comp3360minVal, comp3360minI, comp3360minJ);
    wire [11:0] comp3361minVal;
    wire [5:0] comp3361minI, comp3361minJ;
    Comparator comp3361(comp2996minVal, comp2996minI, comp2996minJ, comp2997minVal, comp2997minI, comp2997minJ, comp3361minVal, comp3361minI, comp3361minJ);
    wire [11:0] comp3362minVal;
    wire [5:0] comp3362minI, comp3362minJ;
    Comparator comp3362(comp2998minVal, comp2998minI, comp2998minJ, comp2999minVal, comp2999minI, comp2999minJ, comp3362minVal, comp3362minI, comp3362minJ);
    wire [11:0] comp3363minVal;
    wire [5:0] comp3363minI, comp3363minJ;
    Comparator comp3363(comp3000minVal, comp3000minI, comp3000minJ, comp3001minVal, comp3001minI, comp3001minJ, comp3363minVal, comp3363minI, comp3363minJ);
    wire [11:0] comp3364minVal;
    wire [5:0] comp3364minI, comp3364minJ;
    Comparator comp3364(comp3002minVal, comp3002minI, comp3002minJ, comp3003minVal, comp3003minI, comp3003minJ, comp3364minVal, comp3364minI, comp3364minJ);
    wire [11:0] comp3365minVal;
    wire [5:0] comp3365minI, comp3365minJ;
    Comparator comp3365(comp3004minVal, comp3004minI, comp3004minJ, comp3005minVal, comp3005minI, comp3005minJ, comp3365minVal, comp3365minI, comp3365minJ);
    wire [11:0] comp3366minVal;
    wire [5:0] comp3366minI, comp3366minJ;
    Comparator comp3366(comp3006minVal, comp3006minI, comp3006minJ, comp3007minVal, comp3007minI, comp3007minJ, comp3366minVal, comp3366minI, comp3366minJ);
    wire [11:0] comp3367minVal;
    wire [5:0] comp3367minI, comp3367minJ;
    Comparator comp3367(comp3008minVal, comp3008minI, comp3008minJ, comp3009minVal, comp3009minI, comp3009minJ, comp3367minVal, comp3367minI, comp3367minJ);
    wire [11:0] comp3368minVal;
    wire [5:0] comp3368minI, comp3368minJ;
    Comparator comp3368(comp3010minVal, comp3010minI, comp3010minJ, comp3011minVal, comp3011minI, comp3011minJ, comp3368minVal, comp3368minI, comp3368minJ);
    wire [11:0] comp3369minVal;
    wire [5:0] comp3369minI, comp3369minJ;
    Comparator comp3369(comp3012minVal, comp3012minI, comp3012minJ, comp3013minVal, comp3013minI, comp3013minJ, comp3369minVal, comp3369minI, comp3369minJ);
    wire [11:0] comp3370minVal;
    wire [5:0] comp3370minI, comp3370minJ;
    Comparator comp3370(comp3014minVal, comp3014minI, comp3014minJ, comp3015minVal, comp3015minI, comp3015minJ, comp3370minVal, comp3370minI, comp3370minJ);
    wire [11:0] comp3371minVal;
    wire [5:0] comp3371minI, comp3371minJ;
    Comparator comp3371(comp3016minVal, comp3016minI, comp3016minJ, comp3017minVal, comp3017minI, comp3017minJ, comp3371minVal, comp3371minI, comp3371minJ);
    wire [11:0] comp3372minVal;
    wire [5:0] comp3372minI, comp3372minJ;
    Comparator comp3372(comp3018minVal, comp3018minI, comp3018minJ, comp3019minVal, comp3019minI, comp3019minJ, comp3372minVal, comp3372minI, comp3372minJ);
    wire [11:0] comp3373minVal;
    wire [5:0] comp3373minI, comp3373minJ;
    Comparator comp3373(comp3020minVal, comp3020minI, comp3020minJ, comp3021minVal, comp3021minI, comp3021minJ, comp3373minVal, comp3373minI, comp3373minJ);
    wire [11:0] comp3374minVal;
    wire [5:0] comp3374minI, comp3374minJ;
    Comparator comp3374(comp3022minVal, comp3022minI, comp3022minJ, comp3023minVal, comp3023minI, comp3023minJ, comp3374minVal, comp3374minI, comp3374minJ);
    wire [11:0] comp3375minVal;
    wire [5:0] comp3375minI, comp3375minJ;
    Comparator comp3375(comp3024minVal, comp3024minI, comp3024minJ, comp3025minVal, comp3025minI, comp3025minJ, comp3375minVal, comp3375minI, comp3375minJ);
    wire [11:0] comp3376minVal;
    wire [5:0] comp3376minI, comp3376minJ;
    Comparator comp3376(comp3026minVal, comp3026minI, comp3026minJ, comp3027minVal, comp3027minI, comp3027minJ, comp3376minVal, comp3376minI, comp3376minJ);
    wire [11:0] comp3377minVal;
    wire [5:0] comp3377minI, comp3377minJ;
    Comparator comp3377(comp3028minVal, comp3028minI, comp3028minJ, comp3029minVal, comp3029minI, comp3029minJ, comp3377minVal, comp3377minI, comp3377minJ);
    wire [11:0] comp3378minVal;
    wire [5:0] comp3378minI, comp3378minJ;
    Comparator comp3378(comp3030minVal, comp3030minI, comp3030minJ, comp3031minVal, comp3031minI, comp3031minJ, comp3378minVal, comp3378minI, comp3378minJ);
    wire [11:0] comp3379minVal;
    wire [5:0] comp3379minI, comp3379minJ;
    Comparator comp3379(comp3032minVal, comp3032minI, comp3032minJ, comp3033minVal, comp3033minI, comp3033minJ, comp3379minVal, comp3379minI, comp3379minJ);
    wire [11:0] comp3380minVal;
    wire [5:0] comp3380minI, comp3380minJ;
    Comparator comp3380(comp3034minVal, comp3034minI, comp3034minJ, comp3035minVal, comp3035minI, comp3035minJ, comp3380minVal, comp3380minI, comp3380minJ);
    wire [11:0] comp3381minVal;
    wire [5:0] comp3381minI, comp3381minJ;
    Comparator comp3381(comp3036minVal, comp3036minI, comp3036minJ, comp3037minVal, comp3037minI, comp3037minJ, comp3381minVal, comp3381minI, comp3381minJ);
    wire [11:0] comp3382minVal;
    wire [5:0] comp3382minI, comp3382minJ;
    Comparator comp3382(comp3038minVal, comp3038minI, comp3038minJ, comp3039minVal, comp3039minI, comp3039minJ, comp3382minVal, comp3382minI, comp3382minJ);
    wire [11:0] comp3383minVal;
    wire [5:0] comp3383minI, comp3383minJ;
    Comparator comp3383(comp3040minVal, comp3040minI, comp3040minJ, comp3041minVal, comp3041minI, comp3041minJ, comp3383minVal, comp3383minI, comp3383minJ);
    wire [11:0] comp3384minVal;
    wire [5:0] comp3384minI, comp3384minJ;
    Comparator comp3384(comp3042minVal, comp3042minI, comp3042minJ, comp3043minVal, comp3043minI, comp3043minJ, comp3384minVal, comp3384minI, comp3384minJ);
    wire [11:0] comp3385minVal;
    wire [5:0] comp3385minI, comp3385minJ;
    Comparator comp3385(comp3044minVal, comp3044minI, comp3044minJ, comp3045minVal, comp3045minI, comp3045minJ, comp3385minVal, comp3385minI, comp3385minJ);
    wire [11:0] comp3386minVal;
    wire [5:0] comp3386minI, comp3386minJ;
    Comparator comp3386(comp3046minVal, comp3046minI, comp3046minJ, comp3047minVal, comp3047minI, comp3047minJ, comp3386minVal, comp3386minI, comp3386minJ);
    wire [11:0] comp3387minVal;
    wire [5:0] comp3387minI, comp3387minJ;
    Comparator comp3387(comp3048minVal, comp3048minI, comp3048minJ, comp3049minVal, comp3049minI, comp3049minJ, comp3387minVal, comp3387minI, comp3387minJ);
    wire [11:0] comp3388minVal;
    wire [5:0] comp3388minI, comp3388minJ;
    Comparator comp3388(comp3050minVal, comp3050minI, comp3050minJ, comp3051minVal, comp3051minI, comp3051minJ, comp3388minVal, comp3388minI, comp3388minJ);
    wire [11:0] comp3389minVal;
    wire [5:0] comp3389minI, comp3389minJ;
    Comparator comp3389(comp3052minVal, comp3052minI, comp3052minJ, comp3053minVal, comp3053minI, comp3053minJ, comp3389minVal, comp3389minI, comp3389minJ);
    wire [11:0] comp3390minVal;
    wire [5:0] comp3390minI, comp3390minJ;
    Comparator comp3390(comp3054minVal, comp3054minI, comp3054minJ, comp3055minVal, comp3055minI, comp3055minJ, comp3390minVal, comp3390minI, comp3390minJ);
    wire [11:0] comp3391minVal;
    wire [5:0] comp3391minI, comp3391minJ;
    Comparator comp3391(comp3056minVal, comp3056minI, comp3056minJ, comp3057minVal, comp3057minI, comp3057minJ, comp3391minVal, comp3391minI, comp3391minJ);
    wire [11:0] comp3392minVal;
    wire [5:0] comp3392minI, comp3392minJ;
    Comparator comp3392(comp3058minVal, comp3058minI, comp3058minJ, comp3059minVal, comp3059minI, comp3059minJ, comp3392minVal, comp3392minI, comp3392minJ);
    wire [11:0] comp3393minVal;
    wire [5:0] comp3393minI, comp3393minJ;
    Comparator comp3393(comp3060minVal, comp3060minI, comp3060minJ, comp3061minVal, comp3061minI, comp3061minJ, comp3393minVal, comp3393minI, comp3393minJ);
    wire [11:0] comp3394minVal;
    wire [5:0] comp3394minI, comp3394minJ;
    Comparator comp3394(comp3062minVal, comp3062minI, comp3062minJ, comp3063minVal, comp3063minI, comp3063minJ, comp3394minVal, comp3394minI, comp3394minJ);
    wire [11:0] comp3395minVal;
    wire [5:0] comp3395minI, comp3395minJ;
    Comparator comp3395(comp3064minVal, comp3064minI, comp3064minJ, comp3065minVal, comp3065minI, comp3065minJ, comp3395minVal, comp3395minI, comp3395minJ);
    wire [11:0] comp3396minVal;
    wire [5:0] comp3396minI, comp3396minJ;
    Comparator comp3396(comp3066minVal, comp3066minI, comp3066minJ, comp3067minVal, comp3067minI, comp3067minJ, comp3396minVal, comp3396minI, comp3396minJ);
    wire [11:0] comp3397minVal;
    wire [5:0] comp3397minI, comp3397minJ;
    Comparator comp3397(comp3068minVal, comp3068minI, comp3068minJ, comp3069minVal, comp3069minI, comp3069minJ, comp3397minVal, comp3397minI, comp3397minJ);
    wire [11:0] comp3398minVal;
    wire [5:0] comp3398minI, comp3398minJ;
    Comparator comp3398(comp3070minVal, comp3070minI, comp3070minJ, comp3071minVal, comp3071minI, comp3071minJ, comp3398minVal, comp3398minI, comp3398minJ);
    wire [11:0] comp3399minVal;
    wire [5:0] comp3399minI, comp3399minJ;
    Comparator comp3399(comp3072minVal, comp3072minI, comp3072minJ, comp3073minVal, comp3073minI, comp3073minJ, comp3399minVal, comp3399minI, comp3399minJ);
    wire [11:0] comp3400minVal;
    wire [5:0] comp3400minI, comp3400minJ;
    Comparator comp3400(comp3074minVal, comp3074minI, comp3074minJ, comp3075minVal, comp3075minI, comp3075minJ, comp3400minVal, comp3400minI, comp3400minJ);
    wire [11:0] comp3401minVal;
    wire [5:0] comp3401minI, comp3401minJ;
    Comparator comp3401(comp3076minVal, comp3076minI, comp3076minJ, comp3077minVal, comp3077minI, comp3077minJ, comp3401minVal, comp3401minI, comp3401minJ);
    wire [11:0] comp3402minVal;
    wire [5:0] comp3402minI, comp3402minJ;
    Comparator comp3402(comp3078minVal, comp3078minI, comp3078minJ, comp3079minVal, comp3079minI, comp3079minJ, comp3402minVal, comp3402minI, comp3402minJ);
    wire [11:0] comp3403minVal;
    wire [5:0] comp3403minI, comp3403minJ;
    Comparator comp3403(comp3080minVal, comp3080minI, comp3080minJ, comp3081minVal, comp3081minI, comp3081minJ, comp3403minVal, comp3403minI, comp3403minJ);
    wire [11:0] comp3404minVal;
    wire [5:0] comp3404minI, comp3404minJ;
    Comparator comp3404(comp3082minVal, comp3082minI, comp3082minJ, comp3083minVal, comp3083minI, comp3083minJ, comp3404minVal, comp3404minI, comp3404minJ);
    wire [11:0] comp3405minVal;
    wire [5:0] comp3405minI, comp3405minJ;
    Comparator comp3405(comp3084minVal, comp3084minI, comp3084minJ, comp3085minVal, comp3085minI, comp3085minJ, comp3405minVal, comp3405minI, comp3405minJ);
    wire [11:0] comp3406minVal;
    wire [5:0] comp3406minI, comp3406minJ;
    Comparator comp3406(comp3086minVal, comp3086minI, comp3086minJ, comp3087minVal, comp3087minI, comp3087minJ, comp3406minVal, comp3406minI, comp3406minJ);
    wire [11:0] comp3407minVal;
    wire [5:0] comp3407minI, comp3407minJ;
    Comparator comp3407(comp3088minVal, comp3088minI, comp3088minJ, comp3089minVal, comp3089minI, comp3089minJ, comp3407minVal, comp3407minI, comp3407minJ);
    wire [11:0] comp3408minVal;
    wire [5:0] comp3408minI, comp3408minJ;
    Comparator comp3408(comp3090minVal, comp3090minI, comp3090minJ, comp3091minVal, comp3091minI, comp3091minJ, comp3408minVal, comp3408minI, comp3408minJ);
    wire [11:0] comp3409minVal;
    wire [5:0] comp3409minI, comp3409minJ;
    Comparator comp3409(comp3092minVal, comp3092minI, comp3092minJ, comp3093minVal, comp3093minI, comp3093minJ, comp3409minVal, comp3409minI, comp3409minJ);
    wire [11:0] comp3410minVal;
    wire [5:0] comp3410minI, comp3410minJ;
    Comparator comp3410(comp3094minVal, comp3094minI, comp3094minJ, comp3095minVal, comp3095minI, comp3095minJ, comp3410minVal, comp3410minI, comp3410minJ);
    wire [11:0] comp3411minVal;
    wire [5:0] comp3411minI, comp3411minJ;
    Comparator comp3411(comp3096minVal, comp3096minI, comp3096minJ, comp3097minVal, comp3097minI, comp3097minJ, comp3411minVal, comp3411minI, comp3411minJ);
    wire [11:0] comp3412minVal;
    wire [5:0] comp3412minI, comp3412minJ;
    Comparator comp3412(comp3098minVal, comp3098minI, comp3098minJ, comp3099minVal, comp3099minI, comp3099minJ, comp3412minVal, comp3412minI, comp3412minJ);
    wire [11:0] comp3413minVal;
    wire [5:0] comp3413minI, comp3413minJ;
    Comparator comp3413(comp3100minVal, comp3100minI, comp3100minJ, comp3101minVal, comp3101minI, comp3101minJ, comp3413minVal, comp3413minI, comp3413minJ);
    wire [11:0] comp3414minVal;
    wire [5:0] comp3414minI, comp3414minJ;
    Comparator comp3414(comp3102minVal, comp3102minI, comp3102minJ, comp3103minVal, comp3103minI, comp3103minJ, comp3414minVal, comp3414minI, comp3414minJ);
    wire [11:0] comp3415minVal;
    wire [5:0] comp3415minI, comp3415minJ;
    Comparator comp3415(comp3104minVal, comp3104minI, comp3104minJ, comp3105minVal, comp3105minI, comp3105minJ, comp3415minVal, comp3415minI, comp3415minJ);
    wire [11:0] comp3416minVal;
    wire [5:0] comp3416minI, comp3416minJ;
    Comparator comp3416(comp3106minVal, comp3106minI, comp3106minJ, comp3107minVal, comp3107minI, comp3107minJ, comp3416minVal, comp3416minI, comp3416minJ);
    wire [11:0] comp3417minVal;
    wire [5:0] comp3417minI, comp3417minJ;
    Comparator comp3417(comp3108minVal, comp3108minI, comp3108minJ, comp3109minVal, comp3109minI, comp3109minJ, comp3417minVal, comp3417minI, comp3417minJ);
    wire [11:0] comp3418minVal;
    wire [5:0] comp3418minI, comp3418minJ;
    Comparator comp3418(comp3110minVal, comp3110minI, comp3110minJ, comp3111minVal, comp3111minI, comp3111minJ, comp3418minVal, comp3418minI, comp3418minJ);
    wire [11:0] comp3419minVal;
    wire [5:0] comp3419minI, comp3419minJ;
    Comparator comp3419(comp3112minVal, comp3112minI, comp3112minJ, comp3113minVal, comp3113minI, comp3113minJ, comp3419minVal, comp3419minI, comp3419minJ);
    wire [11:0] comp3420minVal;
    wire [5:0] comp3420minI, comp3420minJ;
    Comparator comp3420(comp3114minVal, comp3114minI, comp3114minJ, comp3115minVal, comp3115minI, comp3115minJ, comp3420minVal, comp3420minI, comp3420minJ);
    wire [11:0] comp3421minVal;
    wire [5:0] comp3421minI, comp3421minJ;
    Comparator comp3421(comp3116minVal, comp3116minI, comp3116minJ, comp3117minVal, comp3117minI, comp3117minJ, comp3421minVal, comp3421minI, comp3421minJ);
    wire [11:0] comp3422minVal;
    wire [5:0] comp3422minI, comp3422minJ;
    Comparator comp3422(comp3118minVal, comp3118minI, comp3118minJ, comp3119minVal, comp3119minI, comp3119minJ, comp3422minVal, comp3422minI, comp3422minJ);
    wire [11:0] comp3423minVal;
    wire [5:0] comp3423minI, comp3423minJ;
    Comparator comp3423(comp3120minVal, comp3120minI, comp3120minJ, comp3121minVal, comp3121minI, comp3121minJ, comp3423minVal, comp3423minI, comp3423minJ);
    wire [11:0] comp3424minVal;
    wire [5:0] comp3424minI, comp3424minJ;
    Comparator comp3424(comp3122minVal, comp3122minI, comp3122minJ, comp3123minVal, comp3123minI, comp3123minJ, comp3424minVal, comp3424minI, comp3424minJ);
    wire [11:0] comp3425minVal;
    wire [5:0] comp3425minI, comp3425minJ;
    Comparator comp3425(comp3124minVal, comp3124minI, comp3124minJ, comp3125minVal, comp3125minI, comp3125minJ, comp3425minVal, comp3425minI, comp3425minJ);
    wire [11:0] comp3426minVal;
    wire [5:0] comp3426minI, comp3426minJ;
    Comparator comp3426(comp3126minVal, comp3126minI, comp3126minJ, comp3127minVal, comp3127minI, comp3127minJ, comp3426minVal, comp3426minI, comp3426minJ);
    wire [11:0] comp3427minVal;
    wire [5:0] comp3427minI, comp3427minJ;
    Comparator comp3427(comp3128minVal, comp3128minI, comp3128minJ, comp3129minVal, comp3129minI, comp3129minJ, comp3427minVal, comp3427minI, comp3427minJ);
    wire [11:0] comp3428minVal;
    wire [5:0] comp3428minI, comp3428minJ;
    Comparator comp3428(comp3130minVal, comp3130minI, comp3130minJ, comp3131minVal, comp3131minI, comp3131minJ, comp3428minVal, comp3428minI, comp3428minJ);
    wire [11:0] comp3429minVal;
    wire [5:0] comp3429minI, comp3429minJ;
    Comparator comp3429(comp3132minVal, comp3132minI, comp3132minJ, comp3133minVal, comp3133minI, comp3133minJ, comp3429minVal, comp3429minI, comp3429minJ);
    wire [11:0] comp3430minVal;
    wire [5:0] comp3430minI, comp3430minJ;
    Comparator comp3430(comp3134minVal, comp3134minI, comp3134minJ, comp3135minVal, comp3135minI, comp3135minJ, comp3430minVal, comp3430minI, comp3430minJ);
    wire [11:0] comp3431minVal;
    wire [5:0] comp3431minI, comp3431minJ;
    Comparator comp3431(comp3136minVal, comp3136minI, comp3136minJ, comp3137minVal, comp3137minI, comp3137minJ, comp3431minVal, comp3431minI, comp3431minJ);
    wire [11:0] comp3432minVal;
    wire [5:0] comp3432minI, comp3432minJ;
    Comparator comp3432(comp3138minVal, comp3138minI, comp3138minJ, comp3139minVal, comp3139minI, comp3139minJ, comp3432minVal, comp3432minI, comp3432minJ);
    wire [11:0] comp3433minVal;
    wire [5:0] comp3433minI, comp3433minJ;
    Comparator comp3433(comp3140minVal, comp3140minI, comp3140minJ, comp3141minVal, comp3141minI, comp3141minJ, comp3433minVal, comp3433minI, comp3433minJ);
    wire [11:0] comp3434minVal;
    wire [5:0] comp3434minI, comp3434minJ;
    Comparator comp3434(comp3142minVal, comp3142minI, comp3142minJ, comp3143minVal, comp3143minI, comp3143minJ, comp3434minVal, comp3434minI, comp3434minJ);
    wire [11:0] comp3435minVal;
    wire [5:0] comp3435minI, comp3435minJ;
    Comparator comp3435(comp3144minVal, comp3144minI, comp3144minJ, comp3145minVal, comp3145minI, comp3145minJ, comp3435minVal, comp3435minI, comp3435minJ);
    wire [11:0] comp3436minVal;
    wire [5:0] comp3436minI, comp3436minJ;
    Comparator comp3436(comp3146minVal, comp3146minI, comp3146minJ, comp3147minVal, comp3147minI, comp3147minJ, comp3436minVal, comp3436minI, comp3436minJ);
    wire [11:0] comp3437minVal;
    wire [5:0] comp3437minI, comp3437minJ;
    Comparator comp3437(comp3148minVal, comp3148minI, comp3148minJ, comp3149minVal, comp3149minI, comp3149minJ, comp3437minVal, comp3437minI, comp3437minJ);
    wire [11:0] comp3438minVal;
    wire [5:0] comp3438minI, comp3438minJ;
    Comparator comp3438(comp3150minVal, comp3150minI, comp3150minJ, comp3151minVal, comp3151minI, comp3151minJ, comp3438minVal, comp3438minI, comp3438minJ);
    wire [11:0] comp3439minVal;
    wire [5:0] comp3439minI, comp3439minJ;
    Comparator comp3439(comp3152minVal, comp3152minI, comp3152minJ, comp3153minVal, comp3153minI, comp3153minJ, comp3439minVal, comp3439minI, comp3439minJ);
    wire [11:0] comp3440minVal;
    wire [5:0] comp3440minI, comp3440minJ;
    Comparator comp3440(comp3154minVal, comp3154minI, comp3154minJ, comp3155minVal, comp3155minI, comp3155minJ, comp3440minVal, comp3440minI, comp3440minJ);
    wire [11:0] comp3441minVal;
    wire [5:0] comp3441minI, comp3441minJ;
    Comparator comp3441(comp3156minVal, comp3156minI, comp3156minJ, comp3157minVal, comp3157minI, comp3157minJ, comp3441minVal, comp3441minI, comp3441minJ);
    wire [11:0] comp3442minVal;
    wire [5:0] comp3442minI, comp3442minJ;
    Comparator comp3442(comp3158minVal, comp3158minI, comp3158minJ, comp3159minVal, comp3159minI, comp3159minJ, comp3442minVal, comp3442minI, comp3442minJ);
    wire [11:0] comp3443minVal;
    wire [5:0] comp3443minI, comp3443minJ;
    Comparator comp3443(comp3160minVal, comp3160minI, comp3160minJ, comp3161minVal, comp3161minI, comp3161minJ, comp3443minVal, comp3443minI, comp3443minJ);
    wire [11:0] comp3444minVal;
    wire [5:0] comp3444minI, comp3444minJ;
    Comparator comp3444(comp3162minVal, comp3162minI, comp3162minJ, comp3163minVal, comp3163minI, comp3163minJ, comp3444minVal, comp3444minI, comp3444minJ);
    wire [11:0] comp3445minVal;
    wire [5:0] comp3445minI, comp3445minJ;
    Comparator comp3445(comp3164minVal, comp3164minI, comp3164minJ, comp3165minVal, comp3165minI, comp3165minJ, comp3445minVal, comp3445minI, comp3445minJ);
    wire [11:0] comp3446minVal;
    wire [5:0] comp3446minI, comp3446minJ;
    Comparator comp3446(comp3166minVal, comp3166minI, comp3166minJ, comp3167minVal, comp3167minI, comp3167minJ, comp3446minVal, comp3446minI, comp3446minJ);
    wire [11:0] comp3447minVal;
    wire [5:0] comp3447minI, comp3447minJ;
    Comparator comp3447(comp3168minVal, comp3168minI, comp3168minJ, comp3169minVal, comp3169minI, comp3169minJ, comp3447minVal, comp3447minI, comp3447minJ);
    wire [11:0] comp3448minVal;
    wire [5:0] comp3448minI, comp3448minJ;
    Comparator comp3448(comp3170minVal, comp3170minI, comp3170minJ, comp3171minVal, comp3171minI, comp3171minJ, comp3448minVal, comp3448minI, comp3448minJ);
    wire [11:0] comp3449minVal;
    wire [5:0] comp3449minI, comp3449minJ;
    Comparator comp3449(comp3172minVal, comp3172minI, comp3172minJ, comp3173minVal, comp3173minI, comp3173minJ, comp3449minVal, comp3449minI, comp3449minJ);
    wire [11:0] comp3450minVal;
    wire [5:0] comp3450minI, comp3450minJ;
    Comparator comp3450(comp3174minVal, comp3174minI, comp3174minJ, comp3175minVal, comp3175minI, comp3175minJ, comp3450minVal, comp3450minI, comp3450minJ);
    wire [11:0] comp3451minVal;
    wire [5:0] comp3451minI, comp3451minJ;
    Comparator comp3451(comp3176minVal, comp3176minI, comp3176minJ, comp3177minVal, comp3177minI, comp3177minJ, comp3451minVal, comp3451minI, comp3451minJ);
    wire [11:0] comp3452minVal;
    wire [5:0] comp3452minI, comp3452minJ;
    Comparator comp3452(comp3178minVal, comp3178minI, comp3178minJ, comp3179minVal, comp3179minI, comp3179minJ, comp3452minVal, comp3452minI, comp3452minJ);
    wire [11:0] comp3453minVal;
    wire [5:0] comp3453minI, comp3453minJ;
    Comparator comp3453(comp3180minVal, comp3180minI, comp3180minJ, comp3181minVal, comp3181minI, comp3181minJ, comp3453minVal, comp3453minI, comp3453minJ);
    wire [11:0] comp3454minVal;
    wire [5:0] comp3454minI, comp3454minJ;
    Comparator comp3454(comp3182minVal, comp3182minI, comp3182minJ, comp3183minVal, comp3183minI, comp3183minJ, comp3454minVal, comp3454minI, comp3454minJ);
    wire [11:0] comp3455minVal;
    wire [5:0] comp3455minI, comp3455minJ;
    Comparator comp3455(comp3184minVal, comp3184minI, comp3184minJ, comp3185minVal, comp3185minI, comp3185minJ, comp3455minVal, comp3455minI, comp3455minJ);
    wire [11:0] comp3456minVal;
    wire [5:0] comp3456minI, comp3456minJ;
    Comparator comp3456(comp3186minVal, comp3186minI, comp3186minJ, comp3187minVal, comp3187minI, comp3187minJ, comp3456minVal, comp3456minI, comp3456minJ);
    wire [11:0] comp3457minVal;
    wire [5:0] comp3457minI, comp3457minJ;
    Comparator comp3457(comp3188minVal, comp3188minI, comp3188minJ, comp3189minVal, comp3189minI, comp3189minJ, comp3457minVal, comp3457minI, comp3457minJ);
    wire [11:0] comp3458minVal;
    wire [5:0] comp3458minI, comp3458minJ;
    Comparator comp3458(comp3190minVal, comp3190minI, comp3190minJ, comp3191minVal, comp3191minI, comp3191minJ, comp3458minVal, comp3458minI, comp3458minJ);
    wire [11:0] comp3459minVal;
    wire [5:0] comp3459minI, comp3459minJ;
    Comparator comp3459(comp3192minVal, comp3192minI, comp3192minJ, comp3193minVal, comp3193minI, comp3193minJ, comp3459minVal, comp3459minI, comp3459minJ);
    wire [11:0] comp3460minVal;
    wire [5:0] comp3460minI, comp3460minJ;
    Comparator comp3460(comp3194minVal, comp3194minI, comp3194minJ, comp3195minVal, comp3195minI, comp3195minJ, comp3460minVal, comp3460minI, comp3460minJ);
    wire [11:0] comp3461minVal;
    wire [5:0] comp3461minI, comp3461minJ;
    Comparator comp3461(comp3196minVal, comp3196minI, comp3196minJ, comp3197minVal, comp3197minI, comp3197minJ, comp3461minVal, comp3461minI, comp3461minJ);
    wire [11:0] comp3462minVal;
    wire [5:0] comp3462minI, comp3462minJ;
    Comparator comp3462(comp3198minVal, comp3198minI, comp3198minJ, comp3199minVal, comp3199minI, comp3199minJ, comp3462minVal, comp3462minI, comp3462minJ);
    wire [11:0] comp3463minVal;
    wire [5:0] comp3463minI, comp3463minJ;
    Comparator comp3463(comp3200minVal, comp3200minI, comp3200minJ, comp3201minVal, comp3201minI, comp3201minJ, comp3463minVal, comp3463minI, comp3463minJ);
    wire [11:0] comp3464minVal;
    wire [5:0] comp3464minI, comp3464minJ;
    Comparator comp3464(comp3202minVal, comp3202minI, comp3202minJ, comp3203minVal, comp3203minI, comp3203minJ, comp3464minVal, comp3464minI, comp3464minJ);
    wire [11:0] comp3465minVal;
    wire [5:0] comp3465minI, comp3465minJ;
    Comparator comp3465(comp3204minVal, comp3204minI, comp3204minJ, comp3205minVal, comp3205minI, comp3205minJ, comp3465minVal, comp3465minI, comp3465minJ);
    wire [11:0] comp3466minVal;
    wire [5:0] comp3466minI, comp3466minJ;
    Comparator comp3466(comp3206minVal, comp3206minI, comp3206minJ, comp3207minVal, comp3207minI, comp3207minJ, comp3466minVal, comp3466minI, comp3466minJ);
    wire [11:0] comp3467minVal;
    wire [5:0] comp3467minI, comp3467minJ;
    Comparator comp3467(comp3208minVal, comp3208minI, comp3208minJ, comp3209minVal, comp3209minI, comp3209minJ, comp3467minVal, comp3467minI, comp3467minJ);
    wire [11:0] comp3468minVal;
    wire [5:0] comp3468minI, comp3468minJ;
    Comparator comp3468(comp3210minVal, comp3210minI, comp3210minJ, comp3211minVal, comp3211minI, comp3211minJ, comp3468minVal, comp3468minI, comp3468minJ);
    wire [11:0] comp3469minVal;
    wire [5:0] comp3469minI, comp3469minJ;
    Comparator comp3469(comp3212minVal, comp3212minI, comp3212minJ, comp3213minVal, comp3213minI, comp3213minJ, comp3469minVal, comp3469minI, comp3469minJ);
    wire [11:0] comp3470minVal;
    wire [5:0] comp3470minI, comp3470minJ;
    Comparator comp3470(comp3214minVal, comp3214minI, comp3214minJ, comp3215minVal, comp3215minI, comp3215minJ, comp3470minVal, comp3470minI, comp3470minJ);
    wire [11:0] comp3471minVal;
    wire [5:0] comp3471minI, comp3471minJ;
    Comparator comp3471(comp3216minVal, comp3216minI, comp3216minJ, comp3217minVal, comp3217minI, comp3217minJ, comp3471minVal, comp3471minI, comp3471minJ);
    wire [11:0] comp3472minVal;
    wire [5:0] comp3472minI, comp3472minJ;
    Comparator comp3472(comp3218minVal, comp3218minI, comp3218minJ, comp3219minVal, comp3219minI, comp3219minJ, comp3472minVal, comp3472minI, comp3472minJ);
    wire [11:0] comp3473minVal;
    wire [5:0] comp3473minI, comp3473minJ;
    Comparator comp3473(comp3220minVal, comp3220minI, comp3220minJ, comp3221minVal, comp3221minI, comp3221minJ, comp3473minVal, comp3473minI, comp3473minJ);
    wire [11:0] comp3474minVal;
    wire [5:0] comp3474minI, comp3474minJ;
    Comparator comp3474(comp3222minVal, comp3222minI, comp3222minJ, comp3223minVal, comp3223minI, comp3223minJ, comp3474minVal, comp3474minI, comp3474minJ);
    wire [11:0] comp3475minVal;
    wire [5:0] comp3475minI, comp3475minJ;
    Comparator comp3475(comp3224minVal, comp3224minI, comp3224minJ, comp3225minVal, comp3225minI, comp3225minJ, comp3475minVal, comp3475minI, comp3475minJ);
    wire [11:0] comp3476minVal;
    wire [5:0] comp3476minI, comp3476minJ;
    Comparator comp3476(comp3226minVal, comp3226minI, comp3226minJ, comp3227minVal, comp3227minI, comp3227minJ, comp3476minVal, comp3476minI, comp3476minJ);
    wire [11:0] comp3477minVal;
    wire [5:0] comp3477minI, comp3477minJ;
    Comparator comp3477(comp3228minVal, comp3228minI, comp3228minJ, comp3229minVal, comp3229minI, comp3229minJ, comp3477minVal, comp3477minI, comp3477minJ);
    wire [11:0] comp3478minVal;
    wire [5:0] comp3478minI, comp3478minJ;
    Comparator comp3478(comp3230minVal, comp3230minI, comp3230minJ, comp3231minVal, comp3231minI, comp3231minJ, comp3478minVal, comp3478minI, comp3478minJ);
    wire [11:0] comp3479minVal;
    wire [5:0] comp3479minI, comp3479minJ;
    Comparator comp3479(comp3232minVal, comp3232minI, comp3232minJ, comp3233minVal, comp3233minI, comp3233minJ, comp3479minVal, comp3479minI, comp3479minJ);
    wire [11:0] comp3480minVal;
    wire [5:0] comp3480minI, comp3480minJ;
    Comparator comp3480(comp3234minVal, comp3234minI, comp3234minJ, comp3235minVal, comp3235minI, comp3235minJ, comp3480minVal, comp3480minI, comp3480minJ);
    wire [11:0] comp3481minVal;
    wire [5:0] comp3481minI, comp3481minJ;
    Comparator comp3481(comp3236minVal, comp3236minI, comp3236minJ, comp3237minVal, comp3237minI, comp3237minJ, comp3481minVal, comp3481minI, comp3481minJ);
    wire [11:0] comp3482minVal;
    wire [5:0] comp3482minI, comp3482minJ;
    Comparator comp3482(comp3238minVal, comp3238minI, comp3238minJ, comp3239minVal, comp3239minI, comp3239minJ, comp3482minVal, comp3482minI, comp3482minJ);
    wire [11:0] comp3483minVal;
    wire [5:0] comp3483minI, comp3483minJ;
    Comparator comp3483(comp3240minVal, comp3240minI, comp3240minJ, comp3241minVal, comp3241minI, comp3241minJ, comp3483minVal, comp3483minI, comp3483minJ);
    wire [11:0] comp3484minVal;
    wire [5:0] comp3484minI, comp3484minJ;
    Comparator comp3484(comp3242minVal, comp3242minI, comp3242minJ, comp3243minVal, comp3243minI, comp3243minJ, comp3484minVal, comp3484minI, comp3484minJ);
    wire [11:0] comp3485minVal;
    wire [5:0] comp3485minI, comp3485minJ;
    Comparator comp3485(comp3244minVal, comp3244minI, comp3244minJ, comp3245minVal, comp3245minI, comp3245minJ, comp3485minVal, comp3485minI, comp3485minJ);
    wire [11:0] comp3486minVal;
    wire [5:0] comp3486minI, comp3486minJ;
    Comparator comp3486(comp3246minVal, comp3246minI, comp3246minJ, comp3247minVal, comp3247minI, comp3247minJ, comp3486minVal, comp3486minI, comp3486minJ);
    wire [11:0] comp3487minVal;
    wire [5:0] comp3487minI, comp3487minJ;
    Comparator comp3487(comp3248minVal, comp3248minI, comp3248minJ, comp3249minVal, comp3249minI, comp3249minJ, comp3487minVal, comp3487minI, comp3487minJ);
    wire [11:0] comp3488minVal;
    wire [5:0] comp3488minI, comp3488minJ;
    Comparator comp3488(comp3250minVal, comp3250minI, comp3250minJ, comp3251minVal, comp3251minI, comp3251minJ, comp3488minVal, comp3488minI, comp3488minJ);
    wire [11:0] comp3489minVal;
    wire [5:0] comp3489minI, comp3489minJ;
    Comparator comp3489(comp3252minVal, comp3252minI, comp3252minJ, comp3253minVal, comp3253minI, comp3253minJ, comp3489minVal, comp3489minI, comp3489minJ);
    wire [11:0] comp3490minVal;
    wire [5:0] comp3490minI, comp3490minJ;
    Comparator comp3490(comp3254minVal, comp3254minI, comp3254minJ, comp3255minVal, comp3255minI, comp3255minJ, comp3490minVal, comp3490minI, comp3490minJ);
    wire [11:0] comp3491minVal;
    wire [5:0] comp3491minI, comp3491minJ;
    Comparator comp3491(comp3256minVal, comp3256minI, comp3256minJ, comp3257minVal, comp3257minI, comp3257minJ, comp3491minVal, comp3491minI, comp3491minJ);
    wire [11:0] comp3492minVal;
    wire [5:0] comp3492minI, comp3492minJ;
    Comparator comp3492(comp3258minVal, comp3258minI, comp3258minJ, comp3259minVal, comp3259minI, comp3259minJ, comp3492minVal, comp3492minI, comp3492minJ);
    wire [11:0] comp3493minVal;
    wire [5:0] comp3493minI, comp3493minJ;
    assign comp3493minVal = 4095;
    assign comp3493minI = 0;
    assign comp3493minJ = 0;
    wire [11:0] comp3494minVal;
    wire [5:0] comp3494minI, comp3494minJ;
    Comparator comp3494(comp3260minVal, comp3260minI, comp3260minJ, comp3261minVal, comp3261minI, comp3261minJ, comp3494minVal, comp3494minI, comp3494minJ);
    wire [11:0] comp3495minVal;
    wire [5:0] comp3495minI, comp3495minJ;
    Comparator comp3495(comp3262minVal, comp3262minI, comp3262minJ, comp3263minVal, comp3263minI, comp3263minJ, comp3495minVal, comp3495minI, comp3495minJ);
    wire [11:0] comp3496minVal;
    wire [5:0] comp3496minI, comp3496minJ;
    Comparator comp3496(comp3264minVal, comp3264minI, comp3264minJ, comp3265minVal, comp3265minI, comp3265minJ, comp3496minVal, comp3496minI, comp3496minJ);
    wire [11:0] comp3497minVal;
    wire [5:0] comp3497minI, comp3497minJ;
    Comparator comp3497(comp3266minVal, comp3266minI, comp3266minJ, comp3267minVal, comp3267minI, comp3267minJ, comp3497minVal, comp3497minI, comp3497minJ);
    wire [11:0] comp3498minVal;
    wire [5:0] comp3498minI, comp3498minJ;
    Comparator comp3498(comp3268minVal, comp3268minI, comp3268minJ, comp3269minVal, comp3269minI, comp3269minJ, comp3498minVal, comp3498minI, comp3498minJ);
    wire [11:0] comp3499minVal;
    wire [5:0] comp3499minI, comp3499minJ;
    Comparator comp3499(comp3270minVal, comp3270minI, comp3270minJ, comp3271minVal, comp3271minI, comp3271minJ, comp3499minVal, comp3499minI, comp3499minJ);
    wire [11:0] comp3500minVal;
    wire [5:0] comp3500minI, comp3500minJ;
    Comparator comp3500(comp3272minVal, comp3272minI, comp3272minJ, comp3273minVal, comp3273minI, comp3273minJ, comp3500minVal, comp3500minI, comp3500minJ);
    wire [11:0] comp3501minVal;
    wire [5:0] comp3501minI, comp3501minJ;
    Comparator comp3501(comp3274minVal, comp3274minI, comp3274minJ, comp3275minVal, comp3275minI, comp3275minJ, comp3501minVal, comp3501minI, comp3501minJ);
    wire [11:0] comp3502minVal;
    wire [5:0] comp3502minI, comp3502minJ;
    Comparator comp3502(comp3276minVal, comp3276minI, comp3276minJ, comp3277minVal, comp3277minI, comp3277minJ, comp3502minVal, comp3502minI, comp3502minJ);
    wire [11:0] comp3503minVal;
    wire [5:0] comp3503minI, comp3503minJ;
    Comparator comp3503(comp3278minVal, comp3278minI, comp3278minJ, comp3279minVal, comp3279minI, comp3279minJ, comp3503minVal, comp3503minI, comp3503minJ);
    wire [11:0] comp3504minVal;
    wire [5:0] comp3504minI, comp3504minJ;
    Comparator comp3504(comp3280minVal, comp3280minI, comp3280minJ, comp3281minVal, comp3281minI, comp3281minJ, comp3504minVal, comp3504minI, comp3504minJ);
    wire [11:0] comp3505minVal;
    wire [5:0] comp3505minI, comp3505minJ;
    Comparator comp3505(comp3282minVal, comp3282minI, comp3282minJ, comp3283minVal, comp3283minI, comp3283minJ, comp3505minVal, comp3505minI, comp3505minJ);
    wire [11:0] comp3506minVal;
    wire [5:0] comp3506minI, comp3506minJ;
    Comparator comp3506(comp3284minVal, comp3284minI, comp3284minJ, comp3285minVal, comp3285minI, comp3285minJ, comp3506minVal, comp3506minI, comp3506minJ);
    wire [11:0] comp3507minVal;
    wire [5:0] comp3507minI, comp3507minJ;
    Comparator comp3507(comp3286minVal, comp3286minI, comp3286minJ, comp3287minVal, comp3287minI, comp3287minJ, comp3507minVal, comp3507minI, comp3507minJ);
    wire [11:0] comp3508minVal;
    wire [5:0] comp3508minI, comp3508minJ;
    Comparator comp3508(comp3288minVal, comp3288minI, comp3288minJ, comp3289minVal, comp3289minI, comp3289minJ, comp3508minVal, comp3508minI, comp3508minJ);
    wire [11:0] comp3509minVal;
    wire [5:0] comp3509minI, comp3509minJ;
    Comparator comp3509(comp3290minVal, comp3290minI, comp3290minJ, comp3291minVal, comp3291minI, comp3291minJ, comp3509minVal, comp3509minI, comp3509minJ);
    wire [11:0] comp3510minVal;
    wire [5:0] comp3510minI, comp3510minJ;
    Comparator comp3510(comp3292minVal, comp3292minI, comp3292minJ, comp3293minVal, comp3293minI, comp3293minJ, comp3510minVal, comp3510minI, comp3510minJ);
    wire [11:0] comp3511minVal;
    wire [5:0] comp3511minI, comp3511minJ;
    Comparator comp3511(comp3294minVal, comp3294minI, comp3294minJ, comp3295minVal, comp3295minI, comp3295minJ, comp3511minVal, comp3511minI, comp3511minJ);
    wire [11:0] comp3512minVal;
    wire [5:0] comp3512minI, comp3512minJ;
    Comparator comp3512(comp3296minVal, comp3296minI, comp3296minJ, comp3297minVal, comp3297minI, comp3297minJ, comp3512minVal, comp3512minI, comp3512minJ);
    wire [11:0] comp3513minVal;
    wire [5:0] comp3513minI, comp3513minJ;
    Comparator comp3513(comp3298minVal, comp3298minI, comp3298minJ, comp3299minVal, comp3299minI, comp3299minJ, comp3513minVal, comp3513minI, comp3513minJ);
    wire [11:0] comp3514minVal;
    wire [5:0] comp3514minI, comp3514minJ;
    Comparator comp3514(comp3300minVal, comp3300minI, comp3300minJ, comp3301minVal, comp3301minI, comp3301minJ, comp3514minVal, comp3514minI, comp3514minJ);
    wire [11:0] comp3515minVal;
    wire [5:0] comp3515minI, comp3515minJ;
    Comparator comp3515(comp3302minVal, comp3302minI, comp3302minJ, comp3303minVal, comp3303minI, comp3303minJ, comp3515minVal, comp3515minI, comp3515minJ);
    wire [11:0] comp3516minVal;
    wire [5:0] comp3516minI, comp3516minJ;
    Comparator comp3516(comp3304minVal, comp3304minI, comp3304minJ, comp3305minVal, comp3305minI, comp3305minJ, comp3516minVal, comp3516minI, comp3516minJ);
    wire [11:0] comp3517minVal;
    wire [5:0] comp3517minI, comp3517minJ;
    Comparator comp3517(comp3306minVal, comp3306minI, comp3306minJ, comp3307minVal, comp3307minI, comp3307minJ, comp3517minVal, comp3517minI, comp3517minJ);
    wire [11:0] comp3518minVal;
    wire [5:0] comp3518minI, comp3518minJ;
    Comparator comp3518(comp3308minVal, comp3308minI, comp3308minJ, comp3309minVal, comp3309minI, comp3309minJ, comp3518minVal, comp3518minI, comp3518minJ);
    wire [11:0] comp3519minVal;
    wire [5:0] comp3519minI, comp3519minJ;
    Comparator comp3519(comp3310minVal, comp3310minI, comp3310minJ, comp3311minVal, comp3311minI, comp3311minJ, comp3519minVal, comp3519minI, comp3519minJ);
    wire [11:0] comp3520minVal;
    wire [5:0] comp3520minI, comp3520minJ;
    Comparator comp3520(comp3312minVal, comp3312minI, comp3312minJ, comp3313minVal, comp3313minI, comp3313minJ, comp3520minVal, comp3520minI, comp3520minJ);
    wire [11:0] comp3521minVal;
    wire [5:0] comp3521minI, comp3521minJ;
    Comparator comp3521(comp3314minVal, comp3314minI, comp3314minJ, comp3315minVal, comp3315minI, comp3315minJ, comp3521minVal, comp3521minI, comp3521minJ);
    wire [11:0] comp3522minVal;
    wire [5:0] comp3522minI, comp3522minJ;
    Comparator comp3522(comp3316minVal, comp3316minI, comp3316minJ, comp3317minVal, comp3317minI, comp3317minJ, comp3522minVal, comp3522minI, comp3522minJ);
    wire [11:0] comp3523minVal;
    wire [5:0] comp3523minI, comp3523minJ;
    Comparator comp3523(comp3318minVal, comp3318minI, comp3318minJ, comp3319minVal, comp3319minI, comp3319minJ, comp3523minVal, comp3523minI, comp3523minJ);
    wire [11:0] comp3524minVal;
    wire [5:0] comp3524minI, comp3524minJ;
    Comparator comp3524(comp3320minVal, comp3320minI, comp3320minJ, comp3321minVal, comp3321minI, comp3321minJ, comp3524minVal, comp3524minI, comp3524minJ);
    wire [11:0] comp3525minVal;
    wire [5:0] comp3525minI, comp3525minJ;
    Comparator comp3525(comp3322minVal, comp3322minI, comp3322minJ, comp3323minVal, comp3323minI, comp3323minJ, comp3525minVal, comp3525minI, comp3525minJ);
    wire [11:0] comp3526minVal;
    wire [5:0] comp3526minI, comp3526minJ;
    Comparator comp3526(comp3324minVal, comp3324minI, comp3324minJ, comp3325minVal, comp3325minI, comp3325minJ, comp3526minVal, comp3526minI, comp3526minJ);
    wire [11:0] comp3527minVal;
    wire [5:0] comp3527minI, comp3527minJ;
    Comparator comp3527(comp3326minVal, comp3326minI, comp3326minJ, comp3327minVal, comp3327minI, comp3327minJ, comp3527minVal, comp3527minI, comp3527minJ);
    wire [11:0] comp3528minVal;
    wire [5:0] comp3528minI, comp3528minJ;
    Comparator comp3528(comp3328minVal, comp3328minI, comp3328minJ, comp3329minVal, comp3329minI, comp3329minJ, comp3528minVal, comp3528minI, comp3528minJ);
    wire [11:0] comp3529minVal;
    wire [5:0] comp3529minI, comp3529minJ;
    Comparator comp3529(comp3330minVal, comp3330minI, comp3330minJ, comp3331minVal, comp3331minI, comp3331minJ, comp3529minVal, comp3529minI, comp3529minJ);
    wire [11:0] comp3530minVal;
    wire [5:0] comp3530minI, comp3530minJ;
    Comparator comp3530(comp3332minVal, comp3332minI, comp3332minJ, comp3333minVal, comp3333minI, comp3333minJ, comp3530minVal, comp3530minI, comp3530minJ);
    wire [11:0] comp3531minVal;
    wire [5:0] comp3531minI, comp3531minJ;
    Comparator comp3531(comp3334minVal, comp3334minI, comp3334minJ, comp3335minVal, comp3335minI, comp3335minJ, comp3531minVal, comp3531minI, comp3531minJ);
    wire [11:0] comp3532minVal;
    wire [5:0] comp3532minI, comp3532minJ;
    Comparator comp3532(comp3336minVal, comp3336minI, comp3336minJ, comp3337minVal, comp3337minI, comp3337minJ, comp3532minVal, comp3532minI, comp3532minJ);
    wire [11:0] comp3533minVal;
    wire [5:0] comp3533minI, comp3533minJ;
    Comparator comp3533(comp3338minVal, comp3338minI, comp3338minJ, comp3339minVal, comp3339minI, comp3339minJ, comp3533minVal, comp3533minI, comp3533minJ);
    wire [11:0] comp3534minVal;
    wire [5:0] comp3534minI, comp3534minJ;
    Comparator comp3534(comp3340minVal, comp3340minI, comp3340minJ, comp3341minVal, comp3341minI, comp3341minJ, comp3534minVal, comp3534minI, comp3534minJ);
    wire [11:0] comp3535minVal;
    wire [5:0] comp3535minI, comp3535minJ;
    Comparator comp3535(comp3342minVal, comp3342minI, comp3342minJ, comp3343minVal, comp3343minI, comp3343minJ, comp3535minVal, comp3535minI, comp3535minJ);
    wire [11:0] comp3536minVal;
    wire [5:0] comp3536minI, comp3536minJ;
    Comparator comp3536(comp3344minVal, comp3344minI, comp3344minJ, comp3345minVal, comp3345minI, comp3345minJ, comp3536minVal, comp3536minI, comp3536minJ);
    wire [11:0] comp3537minVal;
    wire [5:0] comp3537minI, comp3537minJ;
    Comparator comp3537(comp3346minVal, comp3346minI, comp3346minJ, comp3347minVal, comp3347minI, comp3347minJ, comp3537minVal, comp3537minI, comp3537minJ);
    wire [11:0] comp3538minVal;
    wire [5:0] comp3538minI, comp3538minJ;
    Comparator comp3538(comp3348minVal, comp3348minI, comp3348minJ, comp3349minVal, comp3349minI, comp3349minJ, comp3538minVal, comp3538minI, comp3538minJ);
    wire [11:0] comp3539minVal;
    wire [5:0] comp3539minI, comp3539minJ;
    Comparator comp3539(comp3350minVal, comp3350minI, comp3350minJ, comp3351minVal, comp3351minI, comp3351minJ, comp3539minVal, comp3539minI, comp3539minJ);
    wire [11:0] comp3540minVal;
    wire [5:0] comp3540minI, comp3540minJ;
    Comparator comp3540(comp3352minVal, comp3352minI, comp3352minJ, comp3353minVal, comp3353minI, comp3353minJ, comp3540minVal, comp3540minI, comp3540minJ);
    wire [11:0] comp3541minVal;
    wire [5:0] comp3541minI, comp3541minJ;
    Comparator comp3541(comp3354minVal, comp3354minI, comp3354minJ, comp3355minVal, comp3355minI, comp3355minJ, comp3541minVal, comp3541minI, comp3541minJ);
    wire [11:0] comp3542minVal;
    wire [5:0] comp3542minI, comp3542minJ;
    Comparator comp3542(comp3356minVal, comp3356minI, comp3356minJ, comp3357minVal, comp3357minI, comp3357minJ, comp3542minVal, comp3542minI, comp3542minJ);
    wire [11:0] comp3543minVal;
    wire [5:0] comp3543minI, comp3543minJ;
    Comparator comp3543(comp3358minVal, comp3358minI, comp3358minJ, comp3359minVal, comp3359minI, comp3359minJ, comp3543minVal, comp3543minI, comp3543minJ);
    wire [11:0] comp3544minVal;
    wire [5:0] comp3544minI, comp3544minJ;
    Comparator comp3544(comp3360minVal, comp3360minI, comp3360minJ, comp3361minVal, comp3361minI, comp3361minJ, comp3544minVal, comp3544minI, comp3544minJ);
    wire [11:0] comp3545minVal;
    wire [5:0] comp3545minI, comp3545minJ;
    Comparator comp3545(comp3362minVal, comp3362minI, comp3362minJ, comp3363minVal, comp3363minI, comp3363minJ, comp3545minVal, comp3545minI, comp3545minJ);
    wire [11:0] comp3546minVal;
    wire [5:0] comp3546minI, comp3546minJ;
    Comparator comp3546(comp3364minVal, comp3364minI, comp3364minJ, comp3365minVal, comp3365minI, comp3365minJ, comp3546minVal, comp3546minI, comp3546minJ);
    wire [11:0] comp3547minVal;
    wire [5:0] comp3547minI, comp3547minJ;
    Comparator comp3547(comp3366minVal, comp3366minI, comp3366minJ, comp3367minVal, comp3367minI, comp3367minJ, comp3547minVal, comp3547minI, comp3547minJ);
    wire [11:0] comp3548minVal;
    wire [5:0] comp3548minI, comp3548minJ;
    Comparator comp3548(comp3368minVal, comp3368minI, comp3368minJ, comp3369minVal, comp3369minI, comp3369minJ, comp3548minVal, comp3548minI, comp3548minJ);
    wire [11:0] comp3549minVal;
    wire [5:0] comp3549minI, comp3549minJ;
    Comparator comp3549(comp3370minVal, comp3370minI, comp3370minJ, comp3371minVal, comp3371minI, comp3371minJ, comp3549minVal, comp3549minI, comp3549minJ);
    wire [11:0] comp3550minVal;
    wire [5:0] comp3550minI, comp3550minJ;
    Comparator comp3550(comp3372minVal, comp3372minI, comp3372minJ, comp3373minVal, comp3373minI, comp3373minJ, comp3550minVal, comp3550minI, comp3550minJ);
    wire [11:0] comp3551minVal;
    wire [5:0] comp3551minI, comp3551minJ;
    Comparator comp3551(comp3374minVal, comp3374minI, comp3374minJ, comp3375minVal, comp3375minI, comp3375minJ, comp3551minVal, comp3551minI, comp3551minJ);
    wire [11:0] comp3552minVal;
    wire [5:0] comp3552minI, comp3552minJ;
    Comparator comp3552(comp3376minVal, comp3376minI, comp3376minJ, comp3377minVal, comp3377minI, comp3377minJ, comp3552minVal, comp3552minI, comp3552minJ);
    wire [11:0] comp3553minVal;
    wire [5:0] comp3553minI, comp3553minJ;
    Comparator comp3553(comp3378minVal, comp3378minI, comp3378minJ, comp3379minVal, comp3379minI, comp3379minJ, comp3553minVal, comp3553minI, comp3553minJ);
    wire [11:0] comp3554minVal;
    wire [5:0] comp3554minI, comp3554minJ;
    Comparator comp3554(comp3380minVal, comp3380minI, comp3380minJ, comp3381minVal, comp3381minI, comp3381minJ, comp3554minVal, comp3554minI, comp3554minJ);
    wire [11:0] comp3555minVal;
    wire [5:0] comp3555minI, comp3555minJ;
    Comparator comp3555(comp3382minVal, comp3382minI, comp3382minJ, comp3383minVal, comp3383minI, comp3383minJ, comp3555minVal, comp3555minI, comp3555minJ);
    wire [11:0] comp3556minVal;
    wire [5:0] comp3556minI, comp3556minJ;
    Comparator comp3556(comp3384minVal, comp3384minI, comp3384minJ, comp3385minVal, comp3385minI, comp3385minJ, comp3556minVal, comp3556minI, comp3556minJ);
    wire [11:0] comp3557minVal;
    wire [5:0] comp3557minI, comp3557minJ;
    Comparator comp3557(comp3386minVal, comp3386minI, comp3386minJ, comp3387minVal, comp3387minI, comp3387minJ, comp3557minVal, comp3557minI, comp3557minJ);
    wire [11:0] comp3558minVal;
    wire [5:0] comp3558minI, comp3558minJ;
    Comparator comp3558(comp3388minVal, comp3388minI, comp3388minJ, comp3389minVal, comp3389minI, comp3389minJ, comp3558minVal, comp3558minI, comp3558minJ);
    wire [11:0] comp3559minVal;
    wire [5:0] comp3559minI, comp3559minJ;
    Comparator comp3559(comp3390minVal, comp3390minI, comp3390minJ, comp3391minVal, comp3391minI, comp3391minJ, comp3559minVal, comp3559minI, comp3559minJ);
    wire [11:0] comp3560minVal;
    wire [5:0] comp3560minI, comp3560minJ;
    Comparator comp3560(comp3392minVal, comp3392minI, comp3392minJ, comp3393minVal, comp3393minI, comp3393minJ, comp3560minVal, comp3560minI, comp3560minJ);
    wire [11:0] comp3561minVal;
    wire [5:0] comp3561minI, comp3561minJ;
    Comparator comp3561(comp3394minVal, comp3394minI, comp3394minJ, comp3395minVal, comp3395minI, comp3395minJ, comp3561minVal, comp3561minI, comp3561minJ);
    wire [11:0] comp3562minVal;
    wire [5:0] comp3562minI, comp3562minJ;
    Comparator comp3562(comp3396minVal, comp3396minI, comp3396minJ, comp3397minVal, comp3397minI, comp3397minJ, comp3562minVal, comp3562minI, comp3562minJ);
    wire [11:0] comp3563minVal;
    wire [5:0] comp3563minI, comp3563minJ;
    Comparator comp3563(comp3398minVal, comp3398minI, comp3398minJ, comp3399minVal, comp3399minI, comp3399minJ, comp3563minVal, comp3563minI, comp3563minJ);
    wire [11:0] comp3564minVal;
    wire [5:0] comp3564minI, comp3564minJ;
    Comparator comp3564(comp3400minVal, comp3400minI, comp3400minJ, comp3401minVal, comp3401minI, comp3401minJ, comp3564minVal, comp3564minI, comp3564minJ);
    wire [11:0] comp3565minVal;
    wire [5:0] comp3565minI, comp3565minJ;
    Comparator comp3565(comp3402minVal, comp3402minI, comp3402minJ, comp3403minVal, comp3403minI, comp3403minJ, comp3565minVal, comp3565minI, comp3565minJ);
    wire [11:0] comp3566minVal;
    wire [5:0] comp3566minI, comp3566minJ;
    Comparator comp3566(comp3404minVal, comp3404minI, comp3404minJ, comp3405minVal, comp3405minI, comp3405minJ, comp3566minVal, comp3566minI, comp3566minJ);
    wire [11:0] comp3567minVal;
    wire [5:0] comp3567minI, comp3567minJ;
    Comparator comp3567(comp3406minVal, comp3406minI, comp3406minJ, comp3407minVal, comp3407minI, comp3407minJ, comp3567minVal, comp3567minI, comp3567minJ);
    wire [11:0] comp3568minVal;
    wire [5:0] comp3568minI, comp3568minJ;
    Comparator comp3568(comp3408minVal, comp3408minI, comp3408minJ, comp3409minVal, comp3409minI, comp3409minJ, comp3568minVal, comp3568minI, comp3568minJ);
    wire [11:0] comp3569minVal;
    wire [5:0] comp3569minI, comp3569minJ;
    Comparator comp3569(comp3410minVal, comp3410minI, comp3410minJ, comp3411minVal, comp3411minI, comp3411minJ, comp3569minVal, comp3569minI, comp3569minJ);
    wire [11:0] comp3570minVal;
    wire [5:0] comp3570minI, comp3570minJ;
    Comparator comp3570(comp3412minVal, comp3412minI, comp3412minJ, comp3413minVal, comp3413minI, comp3413minJ, comp3570minVal, comp3570minI, comp3570minJ);
    wire [11:0] comp3571minVal;
    wire [5:0] comp3571minI, comp3571minJ;
    Comparator comp3571(comp3414minVal, comp3414minI, comp3414minJ, comp3415minVal, comp3415minI, comp3415minJ, comp3571minVal, comp3571minI, comp3571minJ);
    wire [11:0] comp3572minVal;
    wire [5:0] comp3572minI, comp3572minJ;
    Comparator comp3572(comp3416minVal, comp3416minI, comp3416minJ, comp3417minVal, comp3417minI, comp3417minJ, comp3572minVal, comp3572minI, comp3572minJ);
    wire [11:0] comp3573minVal;
    wire [5:0] comp3573minI, comp3573minJ;
    Comparator comp3573(comp3418minVal, comp3418minI, comp3418minJ, comp3419minVal, comp3419minI, comp3419minJ, comp3573minVal, comp3573minI, comp3573minJ);
    wire [11:0] comp3574minVal;
    wire [5:0] comp3574minI, comp3574minJ;
    Comparator comp3574(comp3420minVal, comp3420minI, comp3420minJ, comp3421minVal, comp3421minI, comp3421minJ, comp3574minVal, comp3574minI, comp3574minJ);
    wire [11:0] comp3575minVal;
    wire [5:0] comp3575minI, comp3575minJ;
    Comparator comp3575(comp3422minVal, comp3422minI, comp3422minJ, comp3423minVal, comp3423minI, comp3423minJ, comp3575minVal, comp3575minI, comp3575minJ);
    wire [11:0] comp3576minVal;
    wire [5:0] comp3576minI, comp3576minJ;
    Comparator comp3576(comp3424minVal, comp3424minI, comp3424minJ, comp3425minVal, comp3425minI, comp3425minJ, comp3576minVal, comp3576minI, comp3576minJ);
    wire [11:0] comp3577minVal;
    wire [5:0] comp3577minI, comp3577minJ;
    Comparator comp3577(comp3426minVal, comp3426minI, comp3426minJ, comp3427minVal, comp3427minI, comp3427minJ, comp3577minVal, comp3577minI, comp3577minJ);
    wire [11:0] comp3578minVal;
    wire [5:0] comp3578minI, comp3578minJ;
    Comparator comp3578(comp3428minVal, comp3428minI, comp3428minJ, comp3429minVal, comp3429minI, comp3429minJ, comp3578minVal, comp3578minI, comp3578minJ);
    wire [11:0] comp3579minVal;
    wire [5:0] comp3579minI, comp3579minJ;
    Comparator comp3579(comp3430minVal, comp3430minI, comp3430minJ, comp3431minVal, comp3431minI, comp3431minJ, comp3579minVal, comp3579minI, comp3579minJ);
    wire [11:0] comp3580minVal;
    wire [5:0] comp3580minI, comp3580minJ;
    Comparator comp3580(comp3432minVal, comp3432minI, comp3432minJ, comp3433minVal, comp3433minI, comp3433minJ, comp3580minVal, comp3580minI, comp3580minJ);
    wire [11:0] comp3581minVal;
    wire [5:0] comp3581minI, comp3581minJ;
    Comparator comp3581(comp3434minVal, comp3434minI, comp3434minJ, comp3435minVal, comp3435minI, comp3435minJ, comp3581minVal, comp3581minI, comp3581minJ);
    wire [11:0] comp3582minVal;
    wire [5:0] comp3582minI, comp3582minJ;
    Comparator comp3582(comp3436minVal, comp3436minI, comp3436minJ, comp3437minVal, comp3437minI, comp3437minJ, comp3582minVal, comp3582minI, comp3582minJ);
    wire [11:0] comp3583minVal;
    wire [5:0] comp3583minI, comp3583minJ;
    Comparator comp3583(comp3438minVal, comp3438minI, comp3438minJ, comp3439minVal, comp3439minI, comp3439minJ, comp3583minVal, comp3583minI, comp3583minJ);
    wire [11:0] comp3584minVal;
    wire [5:0] comp3584minI, comp3584minJ;
    Comparator comp3584(comp3440minVal, comp3440minI, comp3440minJ, comp3441minVal, comp3441minI, comp3441minJ, comp3584minVal, comp3584minI, comp3584minJ);
    wire [11:0] comp3585minVal;
    wire [5:0] comp3585minI, comp3585minJ;
    Comparator comp3585(comp3442minVal, comp3442minI, comp3442minJ, comp3443minVal, comp3443minI, comp3443minJ, comp3585minVal, comp3585minI, comp3585minJ);
    wire [11:0] comp3586minVal;
    wire [5:0] comp3586minI, comp3586minJ;
    Comparator comp3586(comp3444minVal, comp3444minI, comp3444minJ, comp3445minVal, comp3445minI, comp3445minJ, comp3586minVal, comp3586minI, comp3586minJ);
    wire [11:0] comp3587minVal;
    wire [5:0] comp3587minI, comp3587minJ;
    Comparator comp3587(comp3446minVal, comp3446minI, comp3446minJ, comp3447minVal, comp3447minI, comp3447minJ, comp3587minVal, comp3587minI, comp3587minJ);
    wire [11:0] comp3588minVal;
    wire [5:0] comp3588minI, comp3588minJ;
    Comparator comp3588(comp3448minVal, comp3448minI, comp3448minJ, comp3449minVal, comp3449minI, comp3449minJ, comp3588minVal, comp3588minI, comp3588minJ);
    wire [11:0] comp3589minVal;
    wire [5:0] comp3589minI, comp3589minJ;
    Comparator comp3589(comp3450minVal, comp3450minI, comp3450minJ, comp3451minVal, comp3451minI, comp3451minJ, comp3589minVal, comp3589minI, comp3589minJ);
    wire [11:0] comp3590minVal;
    wire [5:0] comp3590minI, comp3590minJ;
    Comparator comp3590(comp3452minVal, comp3452minI, comp3452minJ, comp3453minVal, comp3453minI, comp3453minJ, comp3590minVal, comp3590minI, comp3590minJ);
    wire [11:0] comp3591minVal;
    wire [5:0] comp3591minI, comp3591minJ;
    Comparator comp3591(comp3454minVal, comp3454minI, comp3454minJ, comp3455minVal, comp3455minI, comp3455minJ, comp3591minVal, comp3591minI, comp3591minJ);
    wire [11:0] comp3592minVal;
    wire [5:0] comp3592minI, comp3592minJ;
    Comparator comp3592(comp3456minVal, comp3456minI, comp3456minJ, comp3457minVal, comp3457minI, comp3457minJ, comp3592minVal, comp3592minI, comp3592minJ);
    wire [11:0] comp3593minVal;
    wire [5:0] comp3593minI, comp3593minJ;
    Comparator comp3593(comp3458minVal, comp3458minI, comp3458minJ, comp3459minVal, comp3459minI, comp3459minJ, comp3593minVal, comp3593minI, comp3593minJ);
    wire [11:0] comp3594minVal;
    wire [5:0] comp3594minI, comp3594minJ;
    Comparator comp3594(comp3460minVal, comp3460minI, comp3460minJ, comp3461minVal, comp3461minI, comp3461minJ, comp3594minVal, comp3594minI, comp3594minJ);
    wire [11:0] comp3595minVal;
    wire [5:0] comp3595minI, comp3595minJ;
    Comparator comp3595(comp3462minVal, comp3462minI, comp3462minJ, comp3463minVal, comp3463minI, comp3463minJ, comp3595minVal, comp3595minI, comp3595minJ);
    wire [11:0] comp3596minVal;
    wire [5:0] comp3596minI, comp3596minJ;
    Comparator comp3596(comp3464minVal, comp3464minI, comp3464minJ, comp3465minVal, comp3465minI, comp3465minJ, comp3596minVal, comp3596minI, comp3596minJ);
    wire [11:0] comp3597minVal;
    wire [5:0] comp3597minI, comp3597minJ;
    Comparator comp3597(comp3466minVal, comp3466minI, comp3466minJ, comp3467minVal, comp3467minI, comp3467minJ, comp3597minVal, comp3597minI, comp3597minJ);
    wire [11:0] comp3598minVal;
    wire [5:0] comp3598minI, comp3598minJ;
    Comparator comp3598(comp3468minVal, comp3468minI, comp3468minJ, comp3469minVal, comp3469minI, comp3469minJ, comp3598minVal, comp3598minI, comp3598minJ);
    wire [11:0] comp3599minVal;
    wire [5:0] comp3599minI, comp3599minJ;
    Comparator comp3599(comp3470minVal, comp3470minI, comp3470minJ, comp3471minVal, comp3471minI, comp3471minJ, comp3599minVal, comp3599minI, comp3599minJ);
    wire [11:0] comp3600minVal;
    wire [5:0] comp3600minI, comp3600minJ;
    Comparator comp3600(comp3472minVal, comp3472minI, comp3472minJ, comp3473minVal, comp3473minI, comp3473minJ, comp3600minVal, comp3600minI, comp3600minJ);
    wire [11:0] comp3601minVal;
    wire [5:0] comp3601minI, comp3601minJ;
    Comparator comp3601(comp3474minVal, comp3474minI, comp3474minJ, comp3475minVal, comp3475minI, comp3475minJ, comp3601minVal, comp3601minI, comp3601minJ);
    wire [11:0] comp3602minVal;
    wire [5:0] comp3602minI, comp3602minJ;
    Comparator comp3602(comp3476minVal, comp3476minI, comp3476minJ, comp3477minVal, comp3477minI, comp3477minJ, comp3602minVal, comp3602minI, comp3602minJ);
    wire [11:0] comp3603minVal;
    wire [5:0] comp3603minI, comp3603minJ;
    Comparator comp3603(comp3478minVal, comp3478minI, comp3478minJ, comp3479minVal, comp3479minI, comp3479minJ, comp3603minVal, comp3603minI, comp3603minJ);
    wire [11:0] comp3604minVal;
    wire [5:0] comp3604minI, comp3604minJ;
    Comparator comp3604(comp3480minVal, comp3480minI, comp3480minJ, comp3481minVal, comp3481minI, comp3481minJ, comp3604minVal, comp3604minI, comp3604minJ);
    wire [11:0] comp3605minVal;
    wire [5:0] comp3605minI, comp3605minJ;
    Comparator comp3605(comp3482minVal, comp3482minI, comp3482minJ, comp3483minVal, comp3483minI, comp3483minJ, comp3605minVal, comp3605minI, comp3605minJ);
    wire [11:0] comp3606minVal;
    wire [5:0] comp3606minI, comp3606minJ;
    Comparator comp3606(comp3484minVal, comp3484minI, comp3484minJ, comp3485minVal, comp3485minI, comp3485minJ, comp3606minVal, comp3606minI, comp3606minJ);
    wire [11:0] comp3607minVal;
    wire [5:0] comp3607minI, comp3607minJ;
    Comparator comp3607(comp3486minVal, comp3486minI, comp3486minJ, comp3487minVal, comp3487minI, comp3487minJ, comp3607minVal, comp3607minI, comp3607minJ);
    wire [11:0] comp3608minVal;
    wire [5:0] comp3608minI, comp3608minJ;
    Comparator comp3608(comp3488minVal, comp3488minI, comp3488minJ, comp3489minVal, comp3489minI, comp3489minJ, comp3608minVal, comp3608minI, comp3608minJ);
    wire [11:0] comp3609minVal;
    wire [5:0] comp3609minI, comp3609minJ;
    Comparator comp3609(comp3490minVal, comp3490minI, comp3490minJ, comp3491minVal, comp3491minI, comp3491minJ, comp3609minVal, comp3609minI, comp3609minJ);
    wire [11:0] comp3610minVal;
    wire [5:0] comp3610minI, comp3610minJ;
    Comparator comp3610(comp3492minVal, comp3492minI, comp3492minJ, comp3493minVal, comp3493minI, comp3493minJ, comp3610minVal, comp3610minI, comp3610minJ);
    wire [11:0] comp3611minVal;
    wire [5:0] comp3611minI, comp3611minJ;
    assign comp3611minVal = 4095;
    assign comp3611minI = 0;
    assign comp3611minJ = 0;
    wire [11:0] comp3612minVal;
    wire [5:0] comp3612minI, comp3612minJ;
    Comparator comp3612(comp3494minVal, comp3494minI, comp3494minJ, comp3495minVal, comp3495minI, comp3495minJ, comp3612minVal, comp3612minI, comp3612minJ);
    wire [11:0] comp3613minVal;
    wire [5:0] comp3613minI, comp3613minJ;
    Comparator comp3613(comp3496minVal, comp3496minI, comp3496minJ, comp3497minVal, comp3497minI, comp3497minJ, comp3613minVal, comp3613minI, comp3613minJ);
    wire [11:0] comp3614minVal;
    wire [5:0] comp3614minI, comp3614minJ;
    Comparator comp3614(comp3498minVal, comp3498minI, comp3498minJ, comp3499minVal, comp3499minI, comp3499minJ, comp3614minVal, comp3614minI, comp3614minJ);
    wire [11:0] comp3615minVal;
    wire [5:0] comp3615minI, comp3615minJ;
    Comparator comp3615(comp3500minVal, comp3500minI, comp3500minJ, comp3501minVal, comp3501minI, comp3501minJ, comp3615minVal, comp3615minI, comp3615minJ);
    wire [11:0] comp3616minVal;
    wire [5:0] comp3616minI, comp3616minJ;
    Comparator comp3616(comp3502minVal, comp3502minI, comp3502minJ, comp3503minVal, comp3503minI, comp3503minJ, comp3616minVal, comp3616minI, comp3616minJ);
    wire [11:0] comp3617minVal;
    wire [5:0] comp3617minI, comp3617minJ;
    Comparator comp3617(comp3504minVal, comp3504minI, comp3504minJ, comp3505minVal, comp3505minI, comp3505minJ, comp3617minVal, comp3617minI, comp3617minJ);
    wire [11:0] comp3618minVal;
    wire [5:0] comp3618minI, comp3618minJ;
    Comparator comp3618(comp3506minVal, comp3506minI, comp3506minJ, comp3507minVal, comp3507minI, comp3507minJ, comp3618minVal, comp3618minI, comp3618minJ);
    wire [11:0] comp3619minVal;
    wire [5:0] comp3619minI, comp3619minJ;
    Comparator comp3619(comp3508minVal, comp3508minI, comp3508minJ, comp3509minVal, comp3509minI, comp3509minJ, comp3619minVal, comp3619minI, comp3619minJ);
    wire [11:0] comp3620minVal;
    wire [5:0] comp3620minI, comp3620minJ;
    Comparator comp3620(comp3510minVal, comp3510minI, comp3510minJ, comp3511minVal, comp3511minI, comp3511minJ, comp3620minVal, comp3620minI, comp3620minJ);
    wire [11:0] comp3621minVal;
    wire [5:0] comp3621minI, comp3621minJ;
    Comparator comp3621(comp3512minVal, comp3512minI, comp3512minJ, comp3513minVal, comp3513minI, comp3513minJ, comp3621minVal, comp3621minI, comp3621minJ);
    wire [11:0] comp3622minVal;
    wire [5:0] comp3622minI, comp3622minJ;
    Comparator comp3622(comp3514minVal, comp3514minI, comp3514minJ, comp3515minVal, comp3515minI, comp3515minJ, comp3622minVal, comp3622minI, comp3622minJ);
    wire [11:0] comp3623minVal;
    wire [5:0] comp3623minI, comp3623minJ;
    Comparator comp3623(comp3516minVal, comp3516minI, comp3516minJ, comp3517minVal, comp3517minI, comp3517minJ, comp3623minVal, comp3623minI, comp3623minJ);
    wire [11:0] comp3624minVal;
    wire [5:0] comp3624minI, comp3624minJ;
    Comparator comp3624(comp3518minVal, comp3518minI, comp3518minJ, comp3519minVal, comp3519minI, comp3519minJ, comp3624minVal, comp3624minI, comp3624minJ);
    wire [11:0] comp3625minVal;
    wire [5:0] comp3625minI, comp3625minJ;
    Comparator comp3625(comp3520minVal, comp3520minI, comp3520minJ, comp3521minVal, comp3521minI, comp3521minJ, comp3625minVal, comp3625minI, comp3625minJ);
    wire [11:0] comp3626minVal;
    wire [5:0] comp3626minI, comp3626minJ;
    Comparator comp3626(comp3522minVal, comp3522minI, comp3522minJ, comp3523minVal, comp3523minI, comp3523minJ, comp3626minVal, comp3626minI, comp3626minJ);
    wire [11:0] comp3627minVal;
    wire [5:0] comp3627minI, comp3627minJ;
    Comparator comp3627(comp3524minVal, comp3524minI, comp3524minJ, comp3525minVal, comp3525minI, comp3525minJ, comp3627minVal, comp3627minI, comp3627minJ);
    wire [11:0] comp3628minVal;
    wire [5:0] comp3628minI, comp3628minJ;
    Comparator comp3628(comp3526minVal, comp3526minI, comp3526minJ, comp3527minVal, comp3527minI, comp3527minJ, comp3628minVal, comp3628minI, comp3628minJ);
    wire [11:0] comp3629minVal;
    wire [5:0] comp3629minI, comp3629minJ;
    Comparator comp3629(comp3528minVal, comp3528minI, comp3528minJ, comp3529minVal, comp3529minI, comp3529minJ, comp3629minVal, comp3629minI, comp3629minJ);
    wire [11:0] comp3630minVal;
    wire [5:0] comp3630minI, comp3630minJ;
    Comparator comp3630(comp3530minVal, comp3530minI, comp3530minJ, comp3531minVal, comp3531minI, comp3531minJ, comp3630minVal, comp3630minI, comp3630minJ);
    wire [11:0] comp3631minVal;
    wire [5:0] comp3631minI, comp3631minJ;
    Comparator comp3631(comp3532minVal, comp3532minI, comp3532minJ, comp3533minVal, comp3533minI, comp3533minJ, comp3631minVal, comp3631minI, comp3631minJ);
    wire [11:0] comp3632minVal;
    wire [5:0] comp3632minI, comp3632minJ;
    Comparator comp3632(comp3534minVal, comp3534minI, comp3534minJ, comp3535minVal, comp3535minI, comp3535minJ, comp3632minVal, comp3632minI, comp3632minJ);
    wire [11:0] comp3633minVal;
    wire [5:0] comp3633minI, comp3633minJ;
    Comparator comp3633(comp3536minVal, comp3536minI, comp3536minJ, comp3537minVal, comp3537minI, comp3537minJ, comp3633minVal, comp3633minI, comp3633minJ);
    wire [11:0] comp3634minVal;
    wire [5:0] comp3634minI, comp3634minJ;
    Comparator comp3634(comp3538minVal, comp3538minI, comp3538minJ, comp3539minVal, comp3539minI, comp3539minJ, comp3634minVal, comp3634minI, comp3634minJ);
    wire [11:0] comp3635minVal;
    wire [5:0] comp3635minI, comp3635minJ;
    Comparator comp3635(comp3540minVal, comp3540minI, comp3540minJ, comp3541minVal, comp3541minI, comp3541minJ, comp3635minVal, comp3635minI, comp3635minJ);
    wire [11:0] comp3636minVal;
    wire [5:0] comp3636minI, comp3636minJ;
    Comparator comp3636(comp3542minVal, comp3542minI, comp3542minJ, comp3543minVal, comp3543minI, comp3543minJ, comp3636minVal, comp3636minI, comp3636minJ);
    wire [11:0] comp3637minVal;
    wire [5:0] comp3637minI, comp3637minJ;
    Comparator comp3637(comp3544minVal, comp3544minI, comp3544minJ, comp3545minVal, comp3545minI, comp3545minJ, comp3637minVal, comp3637minI, comp3637minJ);
    wire [11:0] comp3638minVal;
    wire [5:0] comp3638minI, comp3638minJ;
    Comparator comp3638(comp3546minVal, comp3546minI, comp3546minJ, comp3547minVal, comp3547minI, comp3547minJ, comp3638minVal, comp3638minI, comp3638minJ);
    wire [11:0] comp3639minVal;
    wire [5:0] comp3639minI, comp3639minJ;
    Comparator comp3639(comp3548minVal, comp3548minI, comp3548minJ, comp3549minVal, comp3549minI, comp3549minJ, comp3639minVal, comp3639minI, comp3639minJ);
    wire [11:0] comp3640minVal;
    wire [5:0] comp3640minI, comp3640minJ;
    Comparator comp3640(comp3550minVal, comp3550minI, comp3550minJ, comp3551minVal, comp3551minI, comp3551minJ, comp3640minVal, comp3640minI, comp3640minJ);
    wire [11:0] comp3641minVal;
    wire [5:0] comp3641minI, comp3641minJ;
    Comparator comp3641(comp3552minVal, comp3552minI, comp3552minJ, comp3553minVal, comp3553minI, comp3553minJ, comp3641minVal, comp3641minI, comp3641minJ);
    wire [11:0] comp3642minVal;
    wire [5:0] comp3642minI, comp3642minJ;
    Comparator comp3642(comp3554minVal, comp3554minI, comp3554minJ, comp3555minVal, comp3555minI, comp3555minJ, comp3642minVal, comp3642minI, comp3642minJ);
    wire [11:0] comp3643minVal;
    wire [5:0] comp3643minI, comp3643minJ;
    Comparator comp3643(comp3556minVal, comp3556minI, comp3556minJ, comp3557minVal, comp3557minI, comp3557minJ, comp3643minVal, comp3643minI, comp3643minJ);
    wire [11:0] comp3644minVal;
    wire [5:0] comp3644minI, comp3644minJ;
    Comparator comp3644(comp3558minVal, comp3558minI, comp3558minJ, comp3559minVal, comp3559minI, comp3559minJ, comp3644minVal, comp3644minI, comp3644minJ);
    wire [11:0] comp3645minVal;
    wire [5:0] comp3645minI, comp3645minJ;
    Comparator comp3645(comp3560minVal, comp3560minI, comp3560minJ, comp3561minVal, comp3561minI, comp3561minJ, comp3645minVal, comp3645minI, comp3645minJ);
    wire [11:0] comp3646minVal;
    wire [5:0] comp3646minI, comp3646minJ;
    Comparator comp3646(comp3562minVal, comp3562minI, comp3562minJ, comp3563minVal, comp3563minI, comp3563minJ, comp3646minVal, comp3646minI, comp3646minJ);
    wire [11:0] comp3647minVal;
    wire [5:0] comp3647minI, comp3647minJ;
    Comparator comp3647(comp3564minVal, comp3564minI, comp3564minJ, comp3565minVal, comp3565minI, comp3565minJ, comp3647minVal, comp3647minI, comp3647minJ);
    wire [11:0] comp3648minVal;
    wire [5:0] comp3648minI, comp3648minJ;
    Comparator comp3648(comp3566minVal, comp3566minI, comp3566minJ, comp3567minVal, comp3567minI, comp3567minJ, comp3648minVal, comp3648minI, comp3648minJ);
    wire [11:0] comp3649minVal;
    wire [5:0] comp3649minI, comp3649minJ;
    Comparator comp3649(comp3568minVal, comp3568minI, comp3568minJ, comp3569minVal, comp3569minI, comp3569minJ, comp3649minVal, comp3649minI, comp3649minJ);
    wire [11:0] comp3650minVal;
    wire [5:0] comp3650minI, comp3650minJ;
    Comparator comp3650(comp3570minVal, comp3570minI, comp3570minJ, comp3571minVal, comp3571minI, comp3571minJ, comp3650minVal, comp3650minI, comp3650minJ);
    wire [11:0] comp3651minVal;
    wire [5:0] comp3651minI, comp3651minJ;
    Comparator comp3651(comp3572minVal, comp3572minI, comp3572minJ, comp3573minVal, comp3573minI, comp3573minJ, comp3651minVal, comp3651minI, comp3651minJ);
    wire [11:0] comp3652minVal;
    wire [5:0] comp3652minI, comp3652minJ;
    Comparator comp3652(comp3574minVal, comp3574minI, comp3574minJ, comp3575minVal, comp3575minI, comp3575minJ, comp3652minVal, comp3652minI, comp3652minJ);
    wire [11:0] comp3653minVal;
    wire [5:0] comp3653minI, comp3653minJ;
    Comparator comp3653(comp3576minVal, comp3576minI, comp3576minJ, comp3577minVal, comp3577minI, comp3577minJ, comp3653minVal, comp3653minI, comp3653minJ);
    wire [11:0] comp3654minVal;
    wire [5:0] comp3654minI, comp3654minJ;
    Comparator comp3654(comp3578minVal, comp3578minI, comp3578minJ, comp3579minVal, comp3579minI, comp3579minJ, comp3654minVal, comp3654minI, comp3654minJ);
    wire [11:0] comp3655minVal;
    wire [5:0] comp3655minI, comp3655minJ;
    Comparator comp3655(comp3580minVal, comp3580minI, comp3580minJ, comp3581minVal, comp3581minI, comp3581minJ, comp3655minVal, comp3655minI, comp3655minJ);
    wire [11:0] comp3656minVal;
    wire [5:0] comp3656minI, comp3656minJ;
    Comparator comp3656(comp3582minVal, comp3582minI, comp3582minJ, comp3583minVal, comp3583minI, comp3583minJ, comp3656minVal, comp3656minI, comp3656minJ);
    wire [11:0] comp3657minVal;
    wire [5:0] comp3657minI, comp3657minJ;
    Comparator comp3657(comp3584minVal, comp3584minI, comp3584minJ, comp3585minVal, comp3585minI, comp3585minJ, comp3657minVal, comp3657minI, comp3657minJ);
    wire [11:0] comp3658minVal;
    wire [5:0] comp3658minI, comp3658minJ;
    Comparator comp3658(comp3586minVal, comp3586minI, comp3586minJ, comp3587minVal, comp3587minI, comp3587minJ, comp3658minVal, comp3658minI, comp3658minJ);
    wire [11:0] comp3659minVal;
    wire [5:0] comp3659minI, comp3659minJ;
    Comparator comp3659(comp3588minVal, comp3588minI, comp3588minJ, comp3589minVal, comp3589minI, comp3589minJ, comp3659minVal, comp3659minI, comp3659minJ);
    wire [11:0] comp3660minVal;
    wire [5:0] comp3660minI, comp3660minJ;
    Comparator comp3660(comp3590minVal, comp3590minI, comp3590minJ, comp3591minVal, comp3591minI, comp3591minJ, comp3660minVal, comp3660minI, comp3660minJ);
    wire [11:0] comp3661minVal;
    wire [5:0] comp3661minI, comp3661minJ;
    Comparator comp3661(comp3592minVal, comp3592minI, comp3592minJ, comp3593minVal, comp3593minI, comp3593minJ, comp3661minVal, comp3661minI, comp3661minJ);
    wire [11:0] comp3662minVal;
    wire [5:0] comp3662minI, comp3662minJ;
    Comparator comp3662(comp3594minVal, comp3594minI, comp3594minJ, comp3595minVal, comp3595minI, comp3595minJ, comp3662minVal, comp3662minI, comp3662minJ);
    wire [11:0] comp3663minVal;
    wire [5:0] comp3663minI, comp3663minJ;
    Comparator comp3663(comp3596minVal, comp3596minI, comp3596minJ, comp3597minVal, comp3597minI, comp3597minJ, comp3663minVal, comp3663minI, comp3663minJ);
    wire [11:0] comp3664minVal;
    wire [5:0] comp3664minI, comp3664minJ;
    Comparator comp3664(comp3598minVal, comp3598minI, comp3598minJ, comp3599minVal, comp3599minI, comp3599minJ, comp3664minVal, comp3664minI, comp3664minJ);
    wire [11:0] comp3665minVal;
    wire [5:0] comp3665minI, comp3665minJ;
    Comparator comp3665(comp3600minVal, comp3600minI, comp3600minJ, comp3601minVal, comp3601minI, comp3601minJ, comp3665minVal, comp3665minI, comp3665minJ);
    wire [11:0] comp3666minVal;
    wire [5:0] comp3666minI, comp3666minJ;
    Comparator comp3666(comp3602minVal, comp3602minI, comp3602minJ, comp3603minVal, comp3603minI, comp3603minJ, comp3666minVal, comp3666minI, comp3666minJ);
    wire [11:0] comp3667minVal;
    wire [5:0] comp3667minI, comp3667minJ;
    Comparator comp3667(comp3604minVal, comp3604minI, comp3604minJ, comp3605minVal, comp3605minI, comp3605minJ, comp3667minVal, comp3667minI, comp3667minJ);
    wire [11:0] comp3668minVal;
    wire [5:0] comp3668minI, comp3668minJ;
    Comparator comp3668(comp3606minVal, comp3606minI, comp3606minJ, comp3607minVal, comp3607minI, comp3607minJ, comp3668minVal, comp3668minI, comp3668minJ);
    wire [11:0] comp3669minVal;
    wire [5:0] comp3669minI, comp3669minJ;
    Comparator comp3669(comp3608minVal, comp3608minI, comp3608minJ, comp3609minVal, comp3609minI, comp3609minJ, comp3669minVal, comp3669minI, comp3669minJ);
    wire [11:0] comp3670minVal;
    wire [5:0] comp3670minI, comp3670minJ;
    Comparator comp3670(comp3610minVal, comp3610minI, comp3610minJ, comp3611minVal, comp3611minI, comp3611minJ, comp3670minVal, comp3670minI, comp3670minJ);
    wire [11:0] comp3671minVal;
    wire [5:0] comp3671minI, comp3671minJ;
    assign comp3671minVal = 4095;
    assign comp3671minI = 0;
    assign comp3671minJ = 0;
    wire [11:0] comp3672minVal;
    wire [5:0] comp3672minI, comp3672minJ;
    Comparator comp3672(comp3612minVal, comp3612minI, comp3612minJ, comp3613minVal, comp3613minI, comp3613minJ, comp3672minVal, comp3672minI, comp3672minJ);
    wire [11:0] comp3673minVal;
    wire [5:0] comp3673minI, comp3673minJ;
    Comparator comp3673(comp3614minVal, comp3614minI, comp3614minJ, comp3615minVal, comp3615minI, comp3615minJ, comp3673minVal, comp3673minI, comp3673minJ);
    wire [11:0] comp3674minVal;
    wire [5:0] comp3674minI, comp3674minJ;
    Comparator comp3674(comp3616minVal, comp3616minI, comp3616minJ, comp3617minVal, comp3617minI, comp3617minJ, comp3674minVal, comp3674minI, comp3674minJ);
    wire [11:0] comp3675minVal;
    wire [5:0] comp3675minI, comp3675minJ;
    Comparator comp3675(comp3618minVal, comp3618minI, comp3618minJ, comp3619minVal, comp3619minI, comp3619minJ, comp3675minVal, comp3675minI, comp3675minJ);
    wire [11:0] comp3676minVal;
    wire [5:0] comp3676minI, comp3676minJ;
    Comparator comp3676(comp3620minVal, comp3620minI, comp3620minJ, comp3621minVal, comp3621minI, comp3621minJ, comp3676minVal, comp3676minI, comp3676minJ);
    wire [11:0] comp3677minVal;
    wire [5:0] comp3677minI, comp3677minJ;
    Comparator comp3677(comp3622minVal, comp3622minI, comp3622minJ, comp3623minVal, comp3623minI, comp3623minJ, comp3677minVal, comp3677minI, comp3677minJ);
    wire [11:0] comp3678minVal;
    wire [5:0] comp3678minI, comp3678minJ;
    Comparator comp3678(comp3624minVal, comp3624minI, comp3624minJ, comp3625minVal, comp3625minI, comp3625minJ, comp3678minVal, comp3678minI, comp3678minJ);
    wire [11:0] comp3679minVal;
    wire [5:0] comp3679minI, comp3679minJ;
    Comparator comp3679(comp3626minVal, comp3626minI, comp3626minJ, comp3627minVal, comp3627minI, comp3627minJ, comp3679minVal, comp3679minI, comp3679minJ);
    wire [11:0] comp3680minVal;
    wire [5:0] comp3680minI, comp3680minJ;
    Comparator comp3680(comp3628minVal, comp3628minI, comp3628minJ, comp3629minVal, comp3629minI, comp3629minJ, comp3680minVal, comp3680minI, comp3680minJ);
    wire [11:0] comp3681minVal;
    wire [5:0] comp3681minI, comp3681minJ;
    Comparator comp3681(comp3630minVal, comp3630minI, comp3630minJ, comp3631minVal, comp3631minI, comp3631minJ, comp3681minVal, comp3681minI, comp3681minJ);
    wire [11:0] comp3682minVal;
    wire [5:0] comp3682minI, comp3682minJ;
    Comparator comp3682(comp3632minVal, comp3632minI, comp3632minJ, comp3633minVal, comp3633minI, comp3633minJ, comp3682minVal, comp3682minI, comp3682minJ);
    wire [11:0] comp3683minVal;
    wire [5:0] comp3683minI, comp3683minJ;
    Comparator comp3683(comp3634minVal, comp3634minI, comp3634minJ, comp3635minVal, comp3635minI, comp3635minJ, comp3683minVal, comp3683minI, comp3683minJ);
    wire [11:0] comp3684minVal;
    wire [5:0] comp3684minI, comp3684minJ;
    Comparator comp3684(comp3636minVal, comp3636minI, comp3636minJ, comp3637minVal, comp3637minI, comp3637minJ, comp3684minVal, comp3684minI, comp3684minJ);
    wire [11:0] comp3685minVal;
    wire [5:0] comp3685minI, comp3685minJ;
    Comparator comp3685(comp3638minVal, comp3638minI, comp3638minJ, comp3639minVal, comp3639minI, comp3639minJ, comp3685minVal, comp3685minI, comp3685minJ);
    wire [11:0] comp3686minVal;
    wire [5:0] comp3686minI, comp3686minJ;
    Comparator comp3686(comp3640minVal, comp3640minI, comp3640minJ, comp3641minVal, comp3641minI, comp3641minJ, comp3686minVal, comp3686minI, comp3686minJ);
    wire [11:0] comp3687minVal;
    wire [5:0] comp3687minI, comp3687minJ;
    Comparator comp3687(comp3642minVal, comp3642minI, comp3642minJ, comp3643minVal, comp3643minI, comp3643minJ, comp3687minVal, comp3687minI, comp3687minJ);
    wire [11:0] comp3688minVal;
    wire [5:0] comp3688minI, comp3688minJ;
    Comparator comp3688(comp3644minVal, comp3644minI, comp3644minJ, comp3645minVal, comp3645minI, comp3645minJ, comp3688minVal, comp3688minI, comp3688minJ);
    wire [11:0] comp3689minVal;
    wire [5:0] comp3689minI, comp3689minJ;
    Comparator comp3689(comp3646minVal, comp3646minI, comp3646minJ, comp3647minVal, comp3647minI, comp3647minJ, comp3689minVal, comp3689minI, comp3689minJ);
    wire [11:0] comp3690minVal;
    wire [5:0] comp3690minI, comp3690minJ;
    Comparator comp3690(comp3648minVal, comp3648minI, comp3648minJ, comp3649minVal, comp3649minI, comp3649minJ, comp3690minVal, comp3690minI, comp3690minJ);
    wire [11:0] comp3691minVal;
    wire [5:0] comp3691minI, comp3691minJ;
    Comparator comp3691(comp3650minVal, comp3650minI, comp3650minJ, comp3651minVal, comp3651minI, comp3651minJ, comp3691minVal, comp3691minI, comp3691minJ);
    wire [11:0] comp3692minVal;
    wire [5:0] comp3692minI, comp3692minJ;
    Comparator comp3692(comp3652minVal, comp3652minI, comp3652minJ, comp3653minVal, comp3653minI, comp3653minJ, comp3692minVal, comp3692minI, comp3692minJ);
    wire [11:0] comp3693minVal;
    wire [5:0] comp3693minI, comp3693minJ;
    Comparator comp3693(comp3654minVal, comp3654minI, comp3654minJ, comp3655minVal, comp3655minI, comp3655minJ, comp3693minVal, comp3693minI, comp3693minJ);
    wire [11:0] comp3694minVal;
    wire [5:0] comp3694minI, comp3694minJ;
    Comparator comp3694(comp3656minVal, comp3656minI, comp3656minJ, comp3657minVal, comp3657minI, comp3657minJ, comp3694minVal, comp3694minI, comp3694minJ);
    wire [11:0] comp3695minVal;
    wire [5:0] comp3695minI, comp3695minJ;
    Comparator comp3695(comp3658minVal, comp3658minI, comp3658minJ, comp3659minVal, comp3659minI, comp3659minJ, comp3695minVal, comp3695minI, comp3695minJ);
    wire [11:0] comp3696minVal;
    wire [5:0] comp3696minI, comp3696minJ;
    Comparator comp3696(comp3660minVal, comp3660minI, comp3660minJ, comp3661minVal, comp3661minI, comp3661minJ, comp3696minVal, comp3696minI, comp3696minJ);
    wire [11:0] comp3697minVal;
    wire [5:0] comp3697minI, comp3697minJ;
    Comparator comp3697(comp3662minVal, comp3662minI, comp3662minJ, comp3663minVal, comp3663minI, comp3663minJ, comp3697minVal, comp3697minI, comp3697minJ);
    wire [11:0] comp3698minVal;
    wire [5:0] comp3698minI, comp3698minJ;
    Comparator comp3698(comp3664minVal, comp3664minI, comp3664minJ, comp3665minVal, comp3665minI, comp3665minJ, comp3698minVal, comp3698minI, comp3698minJ);
    wire [11:0] comp3699minVal;
    wire [5:0] comp3699minI, comp3699minJ;
    Comparator comp3699(comp3666minVal, comp3666minI, comp3666minJ, comp3667minVal, comp3667minI, comp3667minJ, comp3699minVal, comp3699minI, comp3699minJ);
    wire [11:0] comp3700minVal;
    wire [5:0] comp3700minI, comp3700minJ;
    Comparator comp3700(comp3668minVal, comp3668minI, comp3668minJ, comp3669minVal, comp3669minI, comp3669minJ, comp3700minVal, comp3700minI, comp3700minJ);
    wire [11:0] comp3701minVal;
    wire [5:0] comp3701minI, comp3701minJ;
    Comparator comp3701(comp3670minVal, comp3670minI, comp3670minJ, comp3671minVal, comp3671minI, comp3671minJ, comp3701minVal, comp3701minI, comp3701minJ);
    wire [11:0] comp3702minVal;
    wire [5:0] comp3702minI, comp3702minJ;
    Comparator comp3702(comp3672minVal, comp3672minI, comp3672minJ, comp3673minVal, comp3673minI, comp3673minJ, comp3702minVal, comp3702minI, comp3702minJ);
    wire [11:0] comp3703minVal;
    wire [5:0] comp3703minI, comp3703minJ;
    Comparator comp3703(comp3674minVal, comp3674minI, comp3674minJ, comp3675minVal, comp3675minI, comp3675minJ, comp3703minVal, comp3703minI, comp3703minJ);
    wire [11:0] comp3704minVal;
    wire [5:0] comp3704minI, comp3704minJ;
    Comparator comp3704(comp3676minVal, comp3676minI, comp3676minJ, comp3677minVal, comp3677minI, comp3677minJ, comp3704minVal, comp3704minI, comp3704minJ);
    wire [11:0] comp3705minVal;
    wire [5:0] comp3705minI, comp3705minJ;
    Comparator comp3705(comp3678minVal, comp3678minI, comp3678minJ, comp3679minVal, comp3679minI, comp3679minJ, comp3705minVal, comp3705minI, comp3705minJ);
    wire [11:0] comp3706minVal;
    wire [5:0] comp3706minI, comp3706minJ;
    Comparator comp3706(comp3680minVal, comp3680minI, comp3680minJ, comp3681minVal, comp3681minI, comp3681minJ, comp3706minVal, comp3706minI, comp3706minJ);
    wire [11:0] comp3707minVal;
    wire [5:0] comp3707minI, comp3707minJ;
    Comparator comp3707(comp3682minVal, comp3682minI, comp3682minJ, comp3683minVal, comp3683minI, comp3683minJ, comp3707minVal, comp3707minI, comp3707minJ);
    wire [11:0] comp3708minVal;
    wire [5:0] comp3708minI, comp3708minJ;
    Comparator comp3708(comp3684minVal, comp3684minI, comp3684minJ, comp3685minVal, comp3685minI, comp3685minJ, comp3708minVal, comp3708minI, comp3708minJ);
    wire [11:0] comp3709minVal;
    wire [5:0] comp3709minI, comp3709minJ;
    Comparator comp3709(comp3686minVal, comp3686minI, comp3686minJ, comp3687minVal, comp3687minI, comp3687minJ, comp3709minVal, comp3709minI, comp3709minJ);
    wire [11:0] comp3710minVal;
    wire [5:0] comp3710minI, comp3710minJ;
    Comparator comp3710(comp3688minVal, comp3688minI, comp3688minJ, comp3689minVal, comp3689minI, comp3689minJ, comp3710minVal, comp3710minI, comp3710minJ);
    wire [11:0] comp3711minVal;
    wire [5:0] comp3711minI, comp3711minJ;
    Comparator comp3711(comp3690minVal, comp3690minI, comp3690minJ, comp3691minVal, comp3691minI, comp3691minJ, comp3711minVal, comp3711minI, comp3711minJ);
    wire [11:0] comp3712minVal;
    wire [5:0] comp3712minI, comp3712minJ;
    Comparator comp3712(comp3692minVal, comp3692minI, comp3692minJ, comp3693minVal, comp3693minI, comp3693minJ, comp3712minVal, comp3712minI, comp3712minJ);
    wire [11:0] comp3713minVal;
    wire [5:0] comp3713minI, comp3713minJ;
    Comparator comp3713(comp3694minVal, comp3694minI, comp3694minJ, comp3695minVal, comp3695minI, comp3695minJ, comp3713minVal, comp3713minI, comp3713minJ);
    wire [11:0] comp3714minVal;
    wire [5:0] comp3714minI, comp3714minJ;
    Comparator comp3714(comp3696minVal, comp3696minI, comp3696minJ, comp3697minVal, comp3697minI, comp3697minJ, comp3714minVal, comp3714minI, comp3714minJ);
    wire [11:0] comp3715minVal;
    wire [5:0] comp3715minI, comp3715minJ;
    Comparator comp3715(comp3698minVal, comp3698minI, comp3698minJ, comp3699minVal, comp3699minI, comp3699minJ, comp3715minVal, comp3715minI, comp3715minJ);
    wire [11:0] comp3716minVal;
    wire [5:0] comp3716minI, comp3716minJ;
    Comparator comp3716(comp3700minVal, comp3700minI, comp3700minJ, comp3701minVal, comp3701minI, comp3701minJ, comp3716minVal, comp3716minI, comp3716minJ);
    wire [11:0] comp3717minVal;
    wire [5:0] comp3717minI, comp3717minJ;
    assign comp3717minVal = 4095;
    assign comp3717minI = 0;
    assign comp3717minJ = 0;
    wire [11:0] comp3718minVal;
    wire [5:0] comp3718minI, comp3718minJ;
    Comparator comp3718(comp3702minVal, comp3702minI, comp3702minJ, comp3703minVal, comp3703minI, comp3703minJ, comp3718minVal, comp3718minI, comp3718minJ);
    wire [11:0] comp3719minVal;
    wire [5:0] comp3719minI, comp3719minJ;
    Comparator comp3719(comp3704minVal, comp3704minI, comp3704minJ, comp3705minVal, comp3705minI, comp3705minJ, comp3719minVal, comp3719minI, comp3719minJ);
    wire [11:0] comp3720minVal;
    wire [5:0] comp3720minI, comp3720minJ;
    Comparator comp3720(comp3706minVal, comp3706minI, comp3706minJ, comp3707minVal, comp3707minI, comp3707minJ, comp3720minVal, comp3720minI, comp3720minJ);
    wire [11:0] comp3721minVal;
    wire [5:0] comp3721minI, comp3721minJ;
    Comparator comp3721(comp3708minVal, comp3708minI, comp3708minJ, comp3709minVal, comp3709minI, comp3709minJ, comp3721minVal, comp3721minI, comp3721minJ);
    wire [11:0] comp3722minVal;
    wire [5:0] comp3722minI, comp3722minJ;
    Comparator comp3722(comp3710minVal, comp3710minI, comp3710minJ, comp3711minVal, comp3711minI, comp3711minJ, comp3722minVal, comp3722minI, comp3722minJ);
    wire [11:0] comp3723minVal;
    wire [5:0] comp3723minI, comp3723minJ;
    Comparator comp3723(comp3712minVal, comp3712minI, comp3712minJ, comp3713minVal, comp3713minI, comp3713minJ, comp3723minVal, comp3723minI, comp3723minJ);
    wire [11:0] comp3724minVal;
    wire [5:0] comp3724minI, comp3724minJ;
    Comparator comp3724(comp3714minVal, comp3714minI, comp3714minJ, comp3715minVal, comp3715minI, comp3715minJ, comp3724minVal, comp3724minI, comp3724minJ);
    wire [11:0] comp3725minVal;
    wire [5:0] comp3725minI, comp3725minJ;
    Comparator comp3725(comp3716minVal, comp3716minI, comp3716minJ, comp3717minVal, comp3717minI, comp3717minJ, comp3725minVal, comp3725minI, comp3725minJ);
    wire [11:0] comp3726minVal;
    wire [5:0] comp3726minI, comp3726minJ;
    Comparator comp3726(comp3718minVal, comp3718minI, comp3718minJ, comp3719minVal, comp3719minI, comp3719minJ, comp3726minVal, comp3726minI, comp3726minJ);
    wire [11:0] comp3727minVal;
    wire [5:0] comp3727minI, comp3727minJ;
    Comparator comp3727(comp3720minVal, comp3720minI, comp3720minJ, comp3721minVal, comp3721minI, comp3721minJ, comp3727minVal, comp3727minI, comp3727minJ);
    wire [11:0] comp3728minVal;
    wire [5:0] comp3728minI, comp3728minJ;
    Comparator comp3728(comp3722minVal, comp3722minI, comp3722minJ, comp3723minVal, comp3723minI, comp3723minJ, comp3728minVal, comp3728minI, comp3728minJ);
    wire [11:0] comp3729minVal;
    wire [5:0] comp3729minI, comp3729minJ;
    Comparator comp3729(comp3724minVal, comp3724minI, comp3724minJ, comp3725minVal, comp3725minI, comp3725minJ, comp3729minVal, comp3729minI, comp3729minJ);
    wire [11:0] comp3730minVal;
    wire [5:0] comp3730minI, comp3730minJ;
    Comparator comp3730(comp3726minVal, comp3726minI, comp3726minJ, comp3727minVal, comp3727minI, comp3727minJ, comp3730minVal, comp3730minI, comp3730minJ);
    wire [11:0] comp3731minVal;
    wire [5:0] comp3731minI, comp3731minJ;
    Comparator comp3731(comp3728minVal, comp3728minI, comp3728minJ, comp3729minVal, comp3729minI, comp3729minJ, comp3731minVal, comp3731minI, comp3731minJ);
    Comparator comp3732(comp3730minVal, comp3730minI, comp3730minJ, comp3731minVal, comp3731minI, comp3731minJ, MinVal, MinI, MinJ);

endmodule
